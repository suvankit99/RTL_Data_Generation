
module square(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] ,
     \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14]
     , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
     \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
     \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
     \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
     \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
     \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
     \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
     \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
     \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
     \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
     \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
     \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
     \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
     \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
     \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
     \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
     \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
     \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
     \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
     \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
     \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
     \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
     \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
     \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
     \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
     \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
     \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
     \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
     \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
     \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
     \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
     \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
     \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103]
     , \asquared[104] , \asquared[105] , \asquared[106] ,
     \asquared[107] , \asquared[108] , \asquared[109] , \asquared[110]
     , \asquared[111] , \asquared[112] , \asquared[113] ,
     \asquared[114] , \asquared[115] , \asquared[116] , \asquared[117]
     , \asquared[118] , \asquared[119] , \asquared[120] ,
     \asquared[121] , \asquared[122] , \asquared[123] , \asquared[124]
     , \asquared[125] , \asquared[126] , \asquared[127] );
  input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
       \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
       \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
       \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
       \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
       \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
       \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
       \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
       \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
       \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
       \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
       \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
       \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
       \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
       \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
       \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
       \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
       \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
       \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
       \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
       \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
       \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
       \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
       \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
       \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
       \asquared[100] , \asquared[101] , \asquared[102] ,
       \asquared[103] , \asquared[104] , \asquared[105] ,
       \asquared[106] , \asquared[107] , \asquared[108] ,
       \asquared[109] , \asquared[110] , \asquared[111] ,
       \asquared[112] , \asquared[113] , \asquared[114] ,
       \asquared[115] , \asquared[116] , \asquared[117] ,
       \asquared[118] , \asquared[119] , \asquared[120] ,
       \asquared[121] , \asquared[122] , \asquared[123] ,
       \asquared[124] , \asquared[125] , \asquared[126] ,
       \asquared[127] ;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  wire \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
       \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
       \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
       \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
       \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
       \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
       \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
       \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
       \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
       \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
       \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
       \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
       \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
       \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
       \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
       \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
       \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
       \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
       \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
       \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
       \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
       \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
       \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
       \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
       \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
       \asquared[100] , \asquared[101] , \asquared[102] ,
       \asquared[103] , \asquared[104] , \asquared[105] ,
       \asquared[106] , \asquared[107] , \asquared[108] ,
       \asquared[109] , \asquared[110] , \asquared[111] ,
       \asquared[112] , \asquared[113] , \asquared[114] ,
       \asquared[115] , \asquared[116] , \asquared[117] ,
       \asquared[118] , \asquared[119] , \asquared[120] ,
       \asquared[121] , \asquared[122] , \asquared[123] ,
       \asquared[124] , \asquared[125] , \asquared[126] ,
       \asquared[127] ;
  wire n194, n196, n197, n198, n200, n201, n202, n203;
  wire n204, n205, n206, n207, n209, n210, n211, n212;
  wire n213, n214, n215, n216, n217, n218, n219, n220;
  wire n221, n223, n224, n225, n226, n227, n228, n229;
  wire n230, n231, n232, n233, n234, n235, n236, n237;
  wire n238, n239, n240, n241, n243, n244, n245, n246;
  wire n247, n248, n249, n250, n251, n252, n253, n254;
  wire n255, n256, n257, n258, n259, n260, n261, n262;
  wire n263, n265, n266, n267, n268, n269, n270, n271;
  wire n272, n273, n274, n275, n276, n277, n278, n279;
  wire n280, n281, n282, n283, n284, n285, n286, n287;
  wire n288, n289, n290, n291, n292, n293, n294, n295;
  wire n296, n298, n299, n300, n301, n302, n303, n304;
  wire n305, n306, n307, n308, n309, n310, n311, n312;
  wire n313, n314, n315, n316, n317, n318, n319, n320;
  wire n321, n322, n323, n324, n325, n326, n327, n328;
  wire n329, n331, n332, n333, n334, n335, n336, n337;
  wire n338, n339, n340, n341, n342, n343, n344, n345;
  wire n346, n347, n348, n349, n350, n351, n352, n353;
  wire n354, n355, n356, n357, n358, n359, n360, n361;
  wire n362, n363, n364, n365, n366, n367, n368, n369;
  wire n370, n371, n372, n373, n375, n376, n377, n378;
  wire n379, n380, n381, n382, n383, n384, n385, n386;
  wire n387, n388, n389, n390, n391, n392, n393, n394;
  wire n395, n396, n397, n398, n399, n400, n401, n402;
  wire n403, n404, n405, n406, n407, n408, n409, n410;
  wire n411, n412, n413, n414, n415, n416, n417, n418;
  wire n419, n421, n422, n423, n424, n425, n426, n427;
  wire n428, n429, n430, n431, n432, n433, n434, n435;
  wire n436, n437, n438, n439, n440, n441, n442, n443;
  wire n444, n445, n446, n447, n448, n449, n450, n451;
  wire n452, n453, n454, n455, n456, n457, n458, n459;
  wire n460, n461, n462, n463, n464, n465, n466, n467;
  wire n468, n469, n470, n471, n473, n474, n475, n476;
  wire n477, n478, n479, n480, n481, n482, n483, n484;
  wire n485, n486, n487, n488, n489, n490, n491, n492;
  wire n493, n494, n495, n496, n497, n498, n499, n500;
  wire n501, n502, n503, n504, n505, n506, n507, n508;
  wire n509, n510, n511, n512, n513, n514, n515, n516;
  wire n517, n518, n519, n520, n521, n522, n523, n524;
  wire n526, n527, n528, n529, n530, n531, n532, n533;
  wire n534, n535, n536, n537, n538, n539, n540, n541;
  wire n542, n543, n544, n545, n546, n547, n548, n549;
  wire n550, n551, n552, n553, n554, n555, n556, n557;
  wire n558, n559, n560, n561, n562, n563, n564, n565;
  wire n566, n567, n568, n569, n570, n571, n572, n573;
  wire n574, n575, n576, n577, n578, n579, n581, n582;
  wire n583, n584, n585, n586, n587, n588, n589, n590;
  wire n591, n592, n593, n594, n595, n596, n597, n598;
  wire n599, n600, n601, n602, n603, n604, n605, n606;
  wire n607, n608, n609, n610, n611, n612, n613, n614;
  wire n615, n616, n617, n618, n619, n620, n621, n622;
  wire n623, n624, n625, n626, n627, n628, n629, n630;
  wire n631, n632, n633, n634, n635, n636, n637, n638;
  wire n639, n640, n641, n642, n643, n644, n646, n647;
  wire n648, n649, n650, n651, n652, n653, n654, n655;
  wire n656, n657, n658, n659, n660, n661, n662, n663;
  wire n664, n667, n668, n669, n670, n671, n672, n673;
  wire n674, n675, n676, n677, n678, n679, n680, n681;
  wire n682, n683, n684, n685, n686, n687, n688, n689;
  wire n690, n691, n692, n693, n694, n695, n696, n697;
  wire n698, n699, n700, n701, n702, n703, n704, n705;
  wire n706, n707, n708, n709, n710, n711, n712, n713;
  wire n714, n716, n717, n718, n719, n720, n721, n722;
  wire n723, n724, n725, n726, n727, n728, n729, n730;
  wire n731, n732, n733, n734, n735, n736, n737, n738;
  wire n739, n740, n741, n742, n743, n744, n745, n746;
  wire n747, n748, n749, n750, n751, n752, n753, n754;
  wire n755, n756, n757, n758, n759, n760, n761, n762;
  wire n763, n764, n765, n766, n767, n768, n769, n770;
  wire n771, n772, n773, n774, n775, n776, n777, n778;
  wire n779, n780, n781, n782, n783, n784, n785, n786;
  wire n787, n788, n789, n791, n792, n793, n794, n795;
  wire n796, n797, n798, n799, n800, n801, n802, n803;
  wire n804, n805, n806, n807, n808, n809, n810, n811;
  wire n812, n813, n814, n815, n816, n817, n818, n819;
  wire n820, n821, n822, n823, n824, n825, n826, n827;
  wire n828, n829, n830, n831, n832, n833, n834, n835;
  wire n836, n837, n838, n839, n840, n841, n842, n843;
  wire n844, n845, n846, n847, n848, n849, n850, n851;
  wire n852, n853, n854, n855, n856, n857, n858, n859;
  wire n860, n861, n862, n863, n864, n865, n866, n867;
  wire n868, n869, n870, n871, n873, n874, n875, n876;
  wire n877, n878, n879, n880, n881, n882, n883, n884;
  wire n885, n886, n887, n888, n889, n890, n891, n892;
  wire n893, n894, n895, n896, n897, n898, n899, n900;
  wire n901, n902, n903, n904, n905, n906, n907, n908;
  wire n909, n910, n911, n912, n913, n914, n915, n916;
  wire n917, n918, n919, n920, n921, n922, n923, n924;
  wire n925, n926, n927, n928, n929, n930, n931, n932;
  wire n933, n934, n935, n936, n937, n938, n939, n940;
  wire n941, n942, n943, n944, n945, n946, n947, n948;
  wire n949, n950, n951, n952, n953, n954, n955, n957;
  wire n958, n959, n960, n961, n962, n963, n964, n965;
  wire n966, n967, n968, n969, n970, n971, n972, n973;
  wire n974, n975, n976, n977, n978, n979, n980, n981;
  wire n982, n983, n984, n985, n986, n987, n988, n989;
  wire n990, n991, n992, n993, n994, n995, n996, n997;
  wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
  wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
  wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  wire n1038, n1039, n1040, n1041, n1042, n1044, n1045, n1046;
  wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
  wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
  wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
  wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
  wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
  wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
  wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
  wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
  wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
  wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
  wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
  wire n1135, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  wire n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151;
  wire n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159;
  wire n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167;
  wire n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175;
  wire n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183;
  wire n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191;
  wire n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199;
  wire n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207;
  wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215;
  wire n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223;
  wire n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231;
  wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
  wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
  wire n1249, n1250, n1251, n1254, n1255, n1256, n1257, n1258;
  wire n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266;
  wire n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274;
  wire n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282;
  wire n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;
  wire n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298;
  wire n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306;
  wire n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314;
  wire n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322;
  wire n1323, n1324, n1325, n1326, n1327, n1329, n1330, n1331;
  wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
  wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
  wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
  wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
  wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
  wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
  wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
  wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
  wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
  wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
  wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
  wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
  wire n1428, n1429, n1431, n1432, n1433, n1434, n1435, n1436;
  wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
  wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
  wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
  wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
  wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
  wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
  wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
  wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
  wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
  wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
  wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
  wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
  wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
  wire n1541, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
  wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
  wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
  wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
  wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
  wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
  wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
  wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
  wire n1606, n1607, n1610, n1611, n1612, n1613, n1614, n1615;
  wire n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623;
  wire n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631;
  wire n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639;
  wire n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647;
  wire n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655;
  wire n1656, n1657, n1658, n1660, n1661, n1662, n1663, n1664;
  wire n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672;
  wire n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680;
  wire n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688;
  wire n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696;
  wire n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704;
  wire n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712;
  wire n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720;
  wire n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728;
  wire n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736;
  wire n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744;
  wire n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752;
  wire n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760;
  wire n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768;
  wire n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776;
  wire n1777, n1778, n1780, n1781, n1782, n1783, n1784, n1785;
  wire n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793;
  wire n1794, n1795, n1796, n1797, n1798, n1799, n1802, n1803;
  wire n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
  wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
  wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827;
  wire n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835;
  wire n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843;
  wire n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
  wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
  wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867;
  wire n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
  wire n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883;
  wire n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891;
  wire n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1900;
  wire n1901, n1902, n1903, n1904, n1905, n1908, n1909, n1910;
  wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
  wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
  wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
  wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
  wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
  wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
  wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
  wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
  wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
  wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
  wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
  wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
  wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
  wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
  wire n2023, n2024, n2026, n2027, n2028, n2029, n2030, n2031;
  wire n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039;
  wire n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047;
  wire n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055;
  wire n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063;
  wire n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071;
  wire n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079;
  wire n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087;
  wire n2088, n2091, n2092, n2093, n2094, n2095, n2096, n2097;
  wire n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105;
  wire n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113;
  wire n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121;
  wire n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129;
  wire n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137;
  wire n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145;
  wire n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153;
  wire n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161;
  wire n2162, n2164, n2165, n2166, n2167, n2168, n2169, n2170;
  wire n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178;
  wire n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186;
  wire n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194;
  wire n2195, n2196, n2197, n2200, n2201, n2202, n2203, n2204;
  wire n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212;
  wire n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220;
  wire n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228;
  wire n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236;
  wire n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244;
  wire n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252;
  wire n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260;
  wire n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268;
  wire n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276;
  wire n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284;
  wire n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292;
  wire n2293, n2294, n2295, n2296, n2298, n2299, n2300, n2301;
  wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
  wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317;
  wire n2318, n2321, n2322, n2323, n2324, n2325, n2326, n2327;
  wire n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335;
  wire n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343;
  wire n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351;
  wire n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359;
  wire n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367;
  wire n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375;
  wire n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383;
  wire n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391;
  wire n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399;
  wire n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407;
  wire n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415;
  wire n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423;
  wire n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431;
  wire n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439;
  wire n2440, n2441, n2442, n2443, n2444, n2446, n2447, n2448;
  wire n2449, n2450, n2451, n2452, n2453, n2454, n2457, n2458;
  wire n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466;
  wire n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474;
  wire n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482;
  wire n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490;
  wire n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498;
  wire n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506;
  wire n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514;
  wire n2515, n2516, n2519, n2520, n2521, n2522, n2523, n2524;
  wire n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532;
  wire n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540;
  wire n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548;
  wire n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556;
  wire n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564;
  wire n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572;
  wire n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580;
  wire n2581, n2582, n2583, n2584, n2586, n2587, n2588, n2589;
  wire n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597;
  wire n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605;
  wire n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613;
  wire n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
  wire n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629;
  wire n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637;
  wire n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645;
  wire n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2655;
  wire n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663;
  wire n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671;
  wire n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679;
  wire n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687;
  wire n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695;
  wire n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703;
  wire n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711;
  wire n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719;
  wire n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727;
  wire n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735;
  wire n2736, n2737, n2738, n2739, n2740, n2742, n2743, n2744;
  wire n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2754;
  wire n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762;
  wire n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770;
  wire n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778;
  wire n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786;
  wire n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794;
  wire n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802;
  wire n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810;
  wire n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818;
  wire n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826;
  wire n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834;
  wire n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842;
  wire n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850;
  wire n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858;
  wire n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866;
  wire n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874;
  wire n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882;
  wire n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890;
  wire n2891, n2892, n2893, n2894, n2895, n2896, n2898, n2899;
  wire n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907;
  wire n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915;
  wire n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923;
  wire n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931;
  wire n2932, n2933, n2934, n2935, n2936, n2939, n2940, n2941;
  wire n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949;
  wire n2950, n2951, n2952, n2955, n2956, n2957, n2958, n2959;
  wire n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967;
  wire n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975;
  wire n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983;
  wire n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991;
  wire n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999;
  wire n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007;
  wire n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015;
  wire n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023;
  wire n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031;
  wire n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039;
  wire n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047;
  wire n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055;
  wire n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064;
  wire n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072;
  wire n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080;
  wire n3081, n3082, n3085, n3086, n3087, n3088, n3089, n3090;
  wire n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098;
  wire n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106;
  wire n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114;
  wire n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122;
  wire n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130;
  wire n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138;
  wire n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146;
  wire n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154;
  wire n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162;
  wire n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170;
  wire n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178;
  wire n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186;
  wire n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194;
  wire n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202;
  wire n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210;
  wire n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218;
  wire n3219, n3220, n3221, n3222, n3224, n3225, n3226, n3227;
  wire n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235;
  wire n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243;
  wire n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251;
  wire n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259;
  wire n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267;
  wire n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275;
  wire n3276, n3277, n3278, n3279, n3280, n3283, n3284, n3285;
  wire n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293;
  wire n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301;
  wire n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309;
  wire n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317;
  wire n3318, n3319, n3320, n3323, n3324, n3325, n3326, n3327;
  wire n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335;
  wire n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343;
  wire n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351;
  wire n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359;
  wire n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367;
  wire n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375;
  wire n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383;
  wire n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391;
  wire n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399;
  wire n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408;
  wire n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416;
  wire n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424;
  wire n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432;
  wire n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440;
  wire n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448;
  wire n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456;
  wire n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464;
  wire n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472;
  wire n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480;
  wire n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488;
  wire n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496;
  wire n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504;
  wire n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512;
  wire n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520;
  wire n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528;
  wire n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536;
  wire n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544;
  wire n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554;
  wire n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562;
  wire n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570;
  wire n3571, n3572, n3573, n3574, n3576, n3577, n3578, n3579;
  wire n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587;
  wire n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595;
  wire n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603;
  wire n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611;
  wire n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619;
  wire n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627;
  wire n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635;
  wire n3636, n3637, n3638, n3639, n3642, n3643, n3644, n3645;
  wire n3646, n3647, n3648, n3649, n3650, n3653, n3654, n3655;
  wire n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663;
  wire n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671;
  wire n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679;
  wire n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687;
  wire n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695;
  wire n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703;
  wire n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711;
  wire n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719;
  wire n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727;
  wire n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735;
  wire n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743;
  wire n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751;
  wire n3752, n3753, n3754, n3755, n3756, n3758, n3759, n3760;
  wire n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768;
  wire n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776;
  wire n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784;
  wire n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792;
  wire n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800;
  wire n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808;
  wire n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816;
  wire n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824;
  wire n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832;
  wire n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840;
  wire n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848;
  wire n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856;
  wire n3857, n3860, n3861, n3862, n3863, n3864, n3865, n3866;
  wire n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874;
  wire n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882;
  wire n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890;
  wire n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898;
  wire n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906;
  wire n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914;
  wire n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922;
  wire n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930;
  wire n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3939;
  wire n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947;
  wire n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955;
  wire n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963;
  wire n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971;
  wire n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979;
  wire n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987;
  wire n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995;
  wire n3996, n3997, n3998, n3999, n4002, n4003, n4004, n4005;
  wire n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013;
  wire n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021;
  wire n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029;
  wire n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037;
  wire n4038, n4041, n4042, n4043, n4044, n4045, n4046, n4047;
  wire n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055;
  wire n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063;
  wire n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071;
  wire n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079;
  wire n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087;
  wire n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095;
  wire n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103;
  wire n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111;
  wire n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119;
  wire n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4128;
  wire n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136;
  wire n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144;
  wire n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152;
  wire n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160;
  wire n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168;
  wire n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176;
  wire n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184;
  wire n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192;
  wire n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200;
  wire n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208;
  wire n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216;
  wire n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224;
  wire n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232;
  wire n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240;
  wire n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248;
  wire n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256;
  wire n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264;
  wire n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272;
  wire n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280;
  wire n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288;
  wire n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296;
  wire n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304;
  wire n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312;
  wire n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320;
  wire n4321, n4322, n4324, n4325, n4326, n4327, n4328, n4329;
  wire n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337;
  wire n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345;
  wire n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353;
  wire n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361;
  wire n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369;
  wire n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377;
  wire n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385;
  wire n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393;
  wire n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401;
  wire n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409;
  wire n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417;
  wire n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425;
  wire n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435;
  wire n4436, n4437, n4438, n4439, n4440, n4441, n4444, n4445;
  wire n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453;
  wire n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461;
  wire n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469;
  wire n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477;
  wire n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485;
  wire n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493;
  wire n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501;
  wire n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509;
  wire n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517;
  wire n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525;
  wire n4526, n4528, n4529, n4530, n4531, n4532, n4533, n4534;
  wire n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544;
  wire n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552;
  wire n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560;
  wire n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568;
  wire n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576;
  wire n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584;
  wire n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592;
  wire n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600;
  wire n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608;
  wire n4609, n4610, n4611, n4612, n4613, n4614, n4617, n4618;
  wire n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626;
  wire n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634;
  wire n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642;
  wire n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650;
  wire n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658;
  wire n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666;
  wire n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674;
  wire n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682;
  wire n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690;
  wire n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698;
  wire n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706;
  wire n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714;
  wire n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722;
  wire n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4731;
  wire n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739;
  wire n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747;
  wire n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755;
  wire n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763;
  wire n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771;
  wire n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779;
  wire n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787;
  wire n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795;
  wire n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803;
  wire n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811;
  wire n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819;
  wire n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827;
  wire n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835;
  wire n4836, n4837, n4838, n4839, n4840, n4841, n4844, n4845;
  wire n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853;
  wire n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861;
  wire n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869;
  wire n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877;
  wire n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885;
  wire n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893;
  wire n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901;
  wire n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909;
  wire n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917;
  wire n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925;
  wire n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933;
  wire n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941;
  wire n4942, n4943, n4944, n4945, n4946, n4947, n4949, n4950;
  wire n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958;
  wire n4959, n4960, n4963, n4964, n4965, n4966, n4967, n4968;
  wire n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976;
  wire n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984;
  wire n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992;
  wire n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000;
  wire n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008;
  wire n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016;
  wire n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024;
  wire n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032;
  wire n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040;
  wire n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048;
  wire n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056;
  wire n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064;
  wire n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072;
  wire n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080;
  wire n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088;
  wire n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096;
  wire n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104;
  wire n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112;
  wire n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120;
  wire n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128;
  wire n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136;
  wire n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144;
  wire n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152;
  wire n5153, n5155, n5156, n5157, n5158, n5159, n5160, n5161;
  wire n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169;
  wire n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177;
  wire n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185;
  wire n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193;
  wire n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201;
  wire n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209;
  wire n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217;
  wire n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225;
  wire n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233;
  wire n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241;
  wire n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249;
  wire n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257;
  wire n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265;
  wire n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273;
  wire n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281;
  wire n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289;
  wire n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297;
  wire n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305;
  wire n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313;
  wire n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321;
  wire n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329;
  wire n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339;
  wire n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347;
  wire n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355;
  wire n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363;
  wire n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371;
  wire n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379;
  wire n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387;
  wire n5388, n5389, n5390, n5392, n5393, n5394, n5395, n5396;
  wire n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404;
  wire n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412;
  wire n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420;
  wire n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428;
  wire n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436;
  wire n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444;
  wire n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452;
  wire n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460;
  wire n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468;
  wire n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476;
  wire n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484;
  wire n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492;
  wire n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500;
  wire n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508;
  wire n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516;
  wire n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524;
  wire n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532;
  wire n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540;
  wire n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548;
  wire n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556;
  wire n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564;
  wire n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572;
  wire n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580;
  wire n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588;
  wire n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596;
  wire n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604;
  wire n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612;
  wire n5613, n5614, n5616, n5617, n5618, n5619, n5620, n5621;
  wire n5622, n5625, n5626, n5627, n5628, n5629, n5630, n5631;
  wire n5632, n5635, n5636, n5637, n5638, n5639, n5640, n5641;
  wire n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649;
  wire n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657;
  wire n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665;
  wire n5666, n5667, n5670, n5671, n5672, n5673, n5674, n5675;
  wire n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683;
  wire n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691;
  wire n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699;
  wire n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707;
  wire n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715;
  wire n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723;
  wire n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731;
  wire n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739;
  wire n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747;
  wire n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755;
  wire n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763;
  wire n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771;
  wire n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779;
  wire n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787;
  wire n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795;
  wire n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803;
  wire n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811;
  wire n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819;
  wire n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827;
  wire n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835;
  wire n5836, n5837, n5838, n5839, n5840, n5842, n5843, n5844;
  wire n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852;
  wire n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860;
  wire n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868;
  wire n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876;
  wire n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884;
  wire n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892;
  wire n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900;
  wire n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908;
  wire n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916;
  wire n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924;
  wire n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932;
  wire n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940;
  wire n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948;
  wire n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956;
  wire n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964;
  wire n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972;
  wire n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980;
  wire n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988;
  wire n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996;
  wire n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004;
  wire n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012;
  wire n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020;
  wire n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028;
  wire n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036;
  wire n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044;
  wire n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052;
  wire n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060;
  wire n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068;
  wire n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6077;
  wire n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085;
  wire n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093;
  wire n6094, n6095, n6096, n6098, n6099, n6100, n6102, n6103;
  wire n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111;
  wire n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119;
  wire n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127;
  wire n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135;
  wire n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143;
  wire n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151;
  wire n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159;
  wire n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167;
  wire n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175;
  wire n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183;
  wire n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191;
  wire n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6201;
  wire n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209;
  wire n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217;
  wire n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225;
  wire n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233;
  wire n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241;
  wire n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249;
  wire n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257;
  wire n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265;
  wire n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273;
  wire n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281;
  wire n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289;
  wire n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297;
  wire n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305;
  wire n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313;
  wire n6314, n6315, n6317, n6318, n6319, n6320, n6321, n6322;
  wire n6323, n6324, n6325, n6326, n6329, n6330, n6331, n6332;
  wire n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340;
  wire n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348;
  wire n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356;
  wire n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364;
  wire n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372;
  wire n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380;
  wire n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388;
  wire n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396;
  wire n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404;
  wire n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412;
  wire n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420;
  wire n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428;
  wire n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436;
  wire n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444;
  wire n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452;
  wire n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460;
  wire n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468;
  wire n6469, n6470, n6471, n6474, n6475, n6476, n6477, n6478;
  wire n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486;
  wire n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494;
  wire n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502;
  wire n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510;
  wire n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518;
  wire n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526;
  wire n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534;
  wire n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542;
  wire n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550;
  wire n6551, n6552, n6553, n6554, n6555, n6557, n6558, n6559;
  wire n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567;
  wire n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575;
  wire n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585;
  wire n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593;
  wire n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601;
  wire n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609;
  wire n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617;
  wire n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625;
  wire n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633;
  wire n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641;
  wire n6642, n6643, n6646, n6647, n6648, n6649, n6650, n6651;
  wire n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659;
  wire n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667;
  wire n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675;
  wire n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683;
  wire n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6693;
  wire n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701;
  wire n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709;
  wire n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717;
  wire n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725;
  wire n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733;
  wire n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741;
  wire n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749;
  wire n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757;
  wire n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765;
  wire n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773;
  wire n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781;
  wire n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789;
  wire n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797;
  wire n6798, n6800, n6801, n6802, n6803, n6804, n6805, n6806;
  wire n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814;
  wire n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822;
  wire n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830;
  wire n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838;
  wire n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846;
  wire n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854;
  wire n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862;
  wire n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870;
  wire n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878;
  wire n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886;
  wire n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894;
  wire n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902;
  wire n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910;
  wire n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918;
  wire n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926;
  wire n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934;
  wire n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942;
  wire n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950;
  wire n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958;
  wire n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966;
  wire n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974;
  wire n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982;
  wire n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990;
  wire n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998;
  wire n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006;
  wire n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014;
  wire n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022;
  wire n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030;
  wire n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038;
  wire n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046;
  wire n7047, n7048, n7049, n7050, n7051, n7052, n7054, n7055;
  wire n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063;
  wire n7064, n7067, n7068, n7069, n7070, n7071, n7072, n7073;
  wire n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081;
  wire n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089;
  wire n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097;
  wire n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105;
  wire n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113;
  wire n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121;
  wire n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129;
  wire n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137;
  wire n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145;
  wire n7146, n7147, n7148, n7151, n7152, n7153, n7154, n7155;
  wire n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163;
  wire n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171;
  wire n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179;
  wire n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187;
  wire n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195;
  wire n7196, n7197, n7198, n7199, n7202, n7203, n7204, n7205;
  wire n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213;
  wire n7214, n7215, n7218, n7219, n7220, n7221, n7222, n7223;
  wire n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231;
  wire n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239;
  wire n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247;
  wire n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255;
  wire n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263;
  wire n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271;
  wire n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279;
  wire n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287;
  wire n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295;
  wire n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303;
  wire n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311;
  wire n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7320;
  wire n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328;
  wire n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336;
  wire n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344;
  wire n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352;
  wire n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360;
  wire n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368;
  wire n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376;
  wire n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384;
  wire n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392;
  wire n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400;
  wire n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408;
  wire n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416;
  wire n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424;
  wire n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432;
  wire n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440;
  wire n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448;
  wire n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456;
  wire n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464;
  wire n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472;
  wire n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480;
  wire n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488;
  wire n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496;
  wire n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504;
  wire n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512;
  wire n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520;
  wire n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528;
  wire n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536;
  wire n7537, n7540, n7541, n7542, n7543, n7544, n7545, n7546;
  wire n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554;
  wire n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562;
  wire n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570;
  wire n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578;
  wire n7579, n7580, n7581, n7582, n7583, n7584, n7586, n7587;
  wire n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595;
  wire n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603;
  wire n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611;
  wire n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619;
  wire n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627;
  wire n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635;
  wire n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643;
  wire n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651;
  wire n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659;
  wire n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667;
  wire n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675;
  wire n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683;
  wire n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691;
  wire n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699;
  wire n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707;
  wire n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715;
  wire n7716, n7719, n7720, n7721, n7722, n7723, n7724, n7725;
  wire n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7735;
  wire n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743;
  wire n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751;
  wire n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759;
  wire n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769;
  wire n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777;
  wire n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785;
  wire n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793;
  wire n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801;
  wire n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809;
  wire n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817;
  wire n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825;
  wire n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833;
  wire n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841;
  wire n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849;
  wire n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857;
  wire n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866;
  wire n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874;
  wire n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882;
  wire n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890;
  wire n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898;
  wire n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906;
  wire n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914;
  wire n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922;
  wire n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930;
  wire n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938;
  wire n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946;
  wire n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954;
  wire n7955, n7956, n7957, n7958, n7959, n7962, n7963, n7964;
  wire n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972;
  wire n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980;
  wire n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988;
  wire n7989, n7990, n7991, n7992, n7993, n7996, n7997, n7998;
  wire n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006;
  wire n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014;
  wire n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022;
  wire n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030;
  wire n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038;
  wire n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046;
  wire n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054;
  wire n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062;
  wire n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070;
  wire n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078;
  wire n8079, n8080, n8081, n8082, n8083, n8084, n8087, n8088;
  wire n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096;
  wire n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104;
  wire n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112;
  wire n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120;
  wire n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129;
  wire n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137;
  wire n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145;
  wire n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153;
  wire n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161;
  wire n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169;
  wire n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177;
  wire n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8187;
  wire n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195;
  wire n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203;
  wire n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211;
  wire n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219;
  wire n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227;
  wire n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235;
  wire n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243;
  wire n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251;
  wire n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259;
  wire n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267;
  wire n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275;
  wire n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283;
  wire n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291;
  wire n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299;
  wire n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307;
  wire n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315;
  wire n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323;
  wire n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331;
  wire n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339;
  wire n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347;
  wire n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355;
  wire n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363;
  wire n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371;
  wire n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379;
  wire n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387;
  wire n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395;
  wire n8396, n8397, n8398, n8399, n8400, n8402, n8403, n8404;
  wire n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412;
  wire n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420;
  wire n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428;
  wire n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436;
  wire n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444;
  wire n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452;
  wire n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460;
  wire n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468;
  wire n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476;
  wire n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484;
  wire n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492;
  wire n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500;
  wire n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508;
  wire n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516;
  wire n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524;
  wire n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532;
  wire n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540;
  wire n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548;
  wire n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556;
  wire n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564;
  wire n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572;
  wire n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580;
  wire n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588;
  wire n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596;
  wire n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604;
  wire n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612;
  wire n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620;
  wire n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628;
  wire n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636;
  wire n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644;
  wire n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652;
  wire n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660;
  wire n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668;
  wire n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676;
  wire n8677, n8678, n8679, n8680, n8681, n8682, n8684, n8685;
  wire n8686, n8687, n8688, n8689, n8690, n8691, n8694, n8695;
  wire n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703;
  wire n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711;
  wire n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719;
  wire n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727;
  wire n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735;
  wire n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743;
  wire n8744, n8745, n8746, n8747, n8748, n8749, n8752, n8753;
  wire n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761;
  wire n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769;
  wire n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777;
  wire n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785;
  wire n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793;
  wire n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801;
  wire n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809;
  wire n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817;
  wire n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825;
  wire n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833;
  wire n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841;
  wire n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849;
  wire n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857;
  wire n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865;
  wire n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873;
  wire n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881;
  wire n8882, n8883, n8884, n8885, n8886, n8889, n8890, n8891;
  wire n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899;
  wire n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907;
  wire n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915;
  wire n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8925;
  wire n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933;
  wire n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941;
  wire n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949;
  wire n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957;
  wire n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965;
  wire n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973;
  wire n8974, n8975, n8977, n8978, n8979, n8980, n8981, n8982;
  wire n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990;
  wire n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998;
  wire n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006;
  wire n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014;
  wire n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022;
  wire n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030;
  wire n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038;
  wire n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046;
  wire n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054;
  wire n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062;
  wire n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070;
  wire n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078;
  wire n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086;
  wire n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094;
  wire n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102;
  wire n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110;
  wire n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118;
  wire n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126;
  wire n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134;
  wire n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142;
  wire n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150;
  wire n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158;
  wire n9159, n9160, n9161, n9162, n9165, n9166, n9167, n9168;
  wire n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176;
  wire n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184;
  wire n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192;
  wire n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200;
  wire n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208;
  wire n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216;
  wire n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224;
  wire n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232;
  wire n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240;
  wire n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248;
  wire n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256;
  wire n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264;
  wire n9265, n9266, n9267, n9268, n9269, n9271, n9272, n9273;
  wire n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281;
  wire n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289;
  wire n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297;
  wire n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305;
  wire n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313;
  wire n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321;
  wire n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329;
  wire n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337;
  wire n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345;
  wire n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353;
  wire n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361;
  wire n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369;
  wire n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377;
  wire n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385;
  wire n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393;
  wire n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401;
  wire n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409;
  wire n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417;
  wire n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425;
  wire n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433;
  wire n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441;
  wire n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449;
  wire n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457;
  wire n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465;
  wire n9466, n9469, n9470, n9471, n9472, n9473, n9474, n9475;
  wire n9476, n9477, n9480, n9481, n9482, n9483, n9484, n9485;
  wire n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493;
  wire n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501;
  wire n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509;
  wire n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517;
  wire n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525;
  wire n9526, n9527, n9528, n9529, n9530, n9533, n9534, n9535;
  wire n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543;
  wire n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551;
  wire n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559;
  wire n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567;
  wire n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576;
  wire n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584;
  wire n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592;
  wire n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600;
  wire n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608;
  wire n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616;
  wire n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624;
  wire n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632;
  wire n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640;
  wire n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648;
  wire n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656;
  wire n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664;
  wire n9665, n9666, n9667, n9670, n9671, n9672, n9673, n9674;
  wire n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682;
  wire n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690;
  wire n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698;
  wire n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706;
  wire n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714;
  wire n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722;
  wire n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730;
  wire n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738;
  wire n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746;
  wire n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754;
  wire n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762;
  wire n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770;
  wire n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778;
  wire n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786;
  wire n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794;
  wire n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802;
  wire n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810;
  wire n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818;
  wire n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826;
  wire n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834;
  wire n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842;
  wire n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850;
  wire n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9859;
  wire n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867;
  wire n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875;
  wire n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883;
  wire n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891;
  wire n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899;
  wire n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907;
  wire n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915;
  wire n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923;
  wire n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931;
  wire n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939;
  wire n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947;
  wire n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955;
  wire n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963;
  wire n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971;
  wire n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979;
  wire n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987;
  wire n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995;
  wire n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003;
  wire n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011;
  wire n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019;
  wire n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027;
  wire n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035;
  wire n10036, n10039, n10040, n10041, n10042, n10043, n10044, n10045;
  wire n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053;
  wire n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061;
  wire n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069;
  wire n10070, n10071, n10072, n10073, n10074, n10075, n10078, n10079;
  wire n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087;
  wire n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095;
  wire n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103;
  wire n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111;
  wire n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119;
  wire n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127;
  wire n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135;
  wire n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143;
  wire n10144, n10145, n10146, n10147, n10149, n10150, n10151, n10152;
  wire n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160;
  wire n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168;
  wire n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176;
  wire n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184;
  wire n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192;
  wire n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200;
  wire n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208;
  wire n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216;
  wire n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224;
  wire n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232;
  wire n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240;
  wire n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248;
  wire n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256;
  wire n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264;
  wire n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272;
  wire n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280;
  wire n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288;
  wire n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296;
  wire n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304;
  wire n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312;
  wire n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320;
  wire n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328;
  wire n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336;
  wire n10337, n10340, n10341, n10342, n10343, n10344, n10345, n10346;
  wire n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10356;
  wire n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364;
  wire n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374;
  wire n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382;
  wire n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390;
  wire n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398;
  wire n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406;
  wire n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414;
  wire n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422;
  wire n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430;
  wire n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439;
  wire n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447;
  wire n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455;
  wire n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463;
  wire n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471;
  wire n10472, n10473, n10474, n10477, n10478, n10479, n10480, n10481;
  wire n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489;
  wire n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497;
  wire n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505;
  wire n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513;
  wire n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521;
  wire n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529;
  wire n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537;
  wire n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545;
  wire n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553;
  wire n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561;
  wire n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569;
  wire n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577;
  wire n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585;
  wire n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593;
  wire n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601;
  wire n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609;
  wire n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617;
  wire n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625;
  wire n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633;
  wire n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641;
  wire n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649;
  wire n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657;
  wire n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665;
  wire n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673;
  wire n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681;
  wire n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689;
  wire n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697;
  wire n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705;
  wire n10706, n10707, n10708, n10709, n10711, n10712, n10713, n10714;
  wire n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722;
  wire n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730;
  wire n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738;
  wire n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746;
  wire n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754;
  wire n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762;
  wire n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770;
  wire n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778;
  wire n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786;
  wire n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794;
  wire n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802;
  wire n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810;
  wire n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818;
  wire n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826;
  wire n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834;
  wire n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842;
  wire n10843, n10844, n10845, n10848, n10849, n10850, n10851, n10852;
  wire n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860;
  wire n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868;
  wire n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876;
  wire n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884;
  wire n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892;
  wire n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900;
  wire n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908;
  wire n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10917;
  wire n10918, n10919, n10921, n10922, n10923, n10924, n10925, n10926;
  wire n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934;
  wire n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942;
  wire n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950;
  wire n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958;
  wire n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966;
  wire n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974;
  wire n10975, n10976, n10978, n10979, n10980, n10981, n10982, n10983;
  wire n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991;
  wire n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999;
  wire n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007;
  wire n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015;
  wire n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023;
  wire n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031;
  wire n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039;
  wire n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047;
  wire n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055;
  wire n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063;
  wire n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071;
  wire n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079;
  wire n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087;
  wire n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095;
  wire n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103;
  wire n11104, n11107, n11108, n11109, n11110, n11111, n11112, n11113;
  wire n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121;
  wire n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129;
  wire n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137;
  wire n11138, n11139, n11140, n11141, n11144, n11145, n11146, n11147;
  wire n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155;
  wire n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163;
  wire n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171;
  wire n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179;
  wire n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187;
  wire n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195;
  wire n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203;
  wire n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211;
  wire n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219;
  wire n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227;
  wire n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235;
  wire n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243;
  wire n11244, n11245, n11246, n11248, n11249, n11250, n11251, n11252;
  wire n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260;
  wire n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268;
  wire n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276;
  wire n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284;
  wire n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292;
  wire n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300;
  wire n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310;
  wire n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318;
  wire n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326;
  wire n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11336;
  wire n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344;
  wire n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352;
  wire n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360;
  wire n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368;
  wire n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376;
  wire n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384;
  wire n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392;
  wire n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400;
  wire n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408;
  wire n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416;
  wire n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424;
  wire n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432;
  wire n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440;
  wire n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448;
  wire n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456;
  wire n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464;
  wire n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472;
  wire n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480;
  wire n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488;
  wire n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496;
  wire n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504;
  wire n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512;
  wire n11513, n11514, n11515, n11517, n11518, n11519, n11520, n11521;
  wire n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529;
  wire n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537;
  wire n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545;
  wire n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553;
  wire n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561;
  wire n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569;
  wire n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577;
  wire n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585;
  wire n11586, n11587, n11588, n11589, n11592, n11593, n11594, n11595;
  wire n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603;
  wire n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611;
  wire n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619;
  wire n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627;
  wire n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635;
  wire n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643;
  wire n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651;
  wire n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659;
  wire n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667;
  wire n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675;
  wire n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683;
  wire n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691;
  wire n11692, n11693, n11694, n11697, n11698, n11699, n11700, n11701;
  wire n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709;
  wire n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717;
  wire n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725;
  wire n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733;
  wire n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741;
  wire n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749;
  wire n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757;
  wire n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765;
  wire n11766, n11767, n11768, n11769, n11771, n11772, n11773, n11774;
  wire n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782;
  wire n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790;
  wire n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798;
  wire n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806;
  wire n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814;
  wire n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822;
  wire n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830;
  wire n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838;
  wire n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846;
  wire n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854;
  wire n11855, n11856, n11857, n11858, n11861, n11862, n11863, n11864;
  wire n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872;
  wire n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880;
  wire n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888;
  wire n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896;
  wire n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904;
  wire n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912;
  wire n11913, n11914, n11917, n11918, n11919, n11920, n11921, n11922;
  wire n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930;
  wire n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938;
  wire n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946;
  wire n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954;
  wire n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962;
  wire n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970;
  wire n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978;
  wire n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986;
  wire n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994;
  wire n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002;
  wire n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010;
  wire n12011, n12012, n12013, n12014, n12015, n12016, n12018, n12019;
  wire n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027;
  wire n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035;
  wire n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043;
  wire n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051;
  wire n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059;
  wire n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067;
  wire n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075;
  wire n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083;
  wire n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091;
  wire n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099;
  wire n12100, n12101, n12102, n12103, n12104, n12107, n12108, n12109;
  wire n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117;
  wire n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125;
  wire n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133;
  wire n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141;
  wire n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149;
  wire n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157;
  wire n12158, n12159, n12160, n12161, n12162, n12163, n12166, n12167;
  wire n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175;
  wire n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183;
  wire n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191;
  wire n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199;
  wire n12200, n12201, n12204, n12205, n12206, n12207, n12208, n12209;
  wire n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217;
  wire n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225;
  wire n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233;
  wire n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241;
  wire n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249;
  wire n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257;
  wire n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12266;
  wire n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274;
  wire n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282;
  wire n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290;
  wire n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298;
  wire n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306;
  wire n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314;
  wire n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322;
  wire n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330;
  wire n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338;
  wire n12339, n12340, n12341, n12342, n12343, n12344, n12347, n12348;
  wire n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356;
  wire n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364;
  wire n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372;
  wire n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380;
  wire n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388;
  wire n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396;
  wire n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404;
  wire n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412;
  wire n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420;
  wire n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428;
  wire n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436;
  wire n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444;
  wire n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452;
  wire n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460;
  wire n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468;
  wire n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476;
  wire n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484;
  wire n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492;
  wire n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500;
  wire n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509;
  wire n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517;
  wire n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525;
  wire n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533;
  wire n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541;
  wire n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12551;
  wire n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559;
  wire n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567;
  wire n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575;
  wire n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583;
  wire n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591;
  wire n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599;
  wire n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607;
  wire n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615;
  wire n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623;
  wire n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631;
  wire n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639;
  wire n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647;
  wire n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655;
  wire n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663;
  wire n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12673;
  wire n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681;
  wire n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689;
  wire n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697;
  wire n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705;
  wire n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713;
  wire n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721;
  wire n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729;
  wire n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737;
  wire n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745;
  wire n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754;
  wire n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762;
  wire n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770;
  wire n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778;
  wire n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786;
  wire n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794;
  wire n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802;
  wire n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810;
  wire n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818;
  wire n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826;
  wire n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834;
  wire n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842;
  wire n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850;
  wire n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858;
  wire n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866;
  wire n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874;
  wire n12875, n12876, n12877, n12878, n12879, n12880, n12883, n12884;
  wire n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892;
  wire n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900;
  wire n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908;
  wire n12909, n12912, n12913, n12914, n12915, n12916, n12917, n12918;
  wire n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926;
  wire n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934;
  wire n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942;
  wire n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950;
  wire n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958;
  wire n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966;
  wire n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974;
  wire n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983;
  wire n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991;
  wire n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999;
  wire n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007;
  wire n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015;
  wire n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023;
  wire n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031;
  wire n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039;
  wire n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047;
  wire n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055;
  wire n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063;
  wire n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071;
  wire n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079;
  wire n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087;
  wire n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095;
  wire n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103;
  wire n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111;
  wire n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119;
  wire n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127;
  wire n13128, n13129, n13130, n13131, n13132, n13135, n13136, n13137;
  wire n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145;
  wire n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153;
  wire n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13163;
  wire n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171;
  wire n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179;
  wire n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187;
  wire n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195;
  wire n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203;
  wire n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212;
  wire n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220;
  wire n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228;
  wire n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236;
  wire n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244;
  wire n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252;
  wire n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260;
  wire n13261, n13262, n13265, n13266, n13267, n13268, n13269, n13270;
  wire n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278;
  wire n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286;
  wire n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294;
  wire n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302;
  wire n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310;
  wire n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318;
  wire n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326;
  wire n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334;
  wire n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342;
  wire n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350;
  wire n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358;
  wire n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366;
  wire n13367, n13368, n13371, n13372, n13373, n13374, n13375, n13376;
  wire n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384;
  wire n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392;
  wire n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400;
  wire n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408;
  wire n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416;
  wire n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424;
  wire n13425, n13426, n13428, n13429, n13430, n13431, n13432, n13433;
  wire n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441;
  wire n13442, n13443, n13444, n13445, n13448, n13449, n13450, n13451;
  wire n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459;
  wire n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467;
  wire n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475;
  wire n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483;
  wire n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491;
  wire n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499;
  wire n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507;
  wire n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515;
  wire n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523;
  wire n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531;
  wire n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539;
  wire n13540, n13541, n13542, n13543, n13544, n13545, n13548, n13549;
  wire n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557;
  wire n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565;
  wire n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573;
  wire n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581;
  wire n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589;
  wire n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597;
  wire n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605;
  wire n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613;
  wire n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621;
  wire n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629;
  wire n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637;
  wire n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645;
  wire n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654;
  wire n13655, n13656, n13657, n13660, n13661, n13662, n13663, n13664;
  wire n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672;
  wire n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680;
  wire n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688;
  wire n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696;
  wire n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704;
  wire n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712;
  wire n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720;
  wire n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728;
  wire n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736;
  wire n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744;
  wire n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752;
  wire n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760;
  wire n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768;
  wire n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776;
  wire n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784;
  wire n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792;
  wire n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800;
  wire n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808;
  wire n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816;
  wire n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824;
  wire n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832;
  wire n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840;
  wire n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848;
  wire n13849, n13850, n13851, n13852, n13853, n13854, n13856, n13857;
  wire n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865;
  wire n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873;
  wire n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881;
  wire n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889;
  wire n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897;
  wire n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905;
  wire n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913;
  wire n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921;
  wire n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929;
  wire n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937;
  wire n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945;
  wire n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953;
  wire n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961;
  wire n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969;
  wire n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977;
  wire n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985;
  wire n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993;
  wire n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001;
  wire n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009;
  wire n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017;
  wire n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025;
  wire n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033;
  wire n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041;
  wire n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049;
  wire n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057;
  wire n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065;
  wire n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14074;
  wire n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082;
  wire n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090;
  wire n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098;
  wire n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106;
  wire n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114;
  wire n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122;
  wire n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130;
  wire n14131, n14132, n14133, n14134, n14135, n14138, n14139, n14140;
  wire n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148;
  wire n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156;
  wire n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164;
  wire n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172;
  wire n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180;
  wire n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188;
  wire n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196;
  wire n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204;
  wire n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212;
  wire n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220;
  wire n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228;
  wire n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236;
  wire n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244;
  wire n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252;
  wire n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260;
  wire n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268;
  wire n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276;
  wire n14277, n14279, n14280, n14281, n14282, n14283, n14284, n14285;
  wire n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293;
  wire n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301;
  wire n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309;
  wire n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317;
  wire n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325;
  wire n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333;
  wire n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341;
  wire n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349;
  wire n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357;
  wire n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365;
  wire n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373;
  wire n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14383;
  wire n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391;
  wire n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399;
  wire n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407;
  wire n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415;
  wire n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423;
  wire n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431;
  wire n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439;
  wire n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447;
  wire n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455;
  wire n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463;
  wire n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471;
  wire n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479;
  wire n14480, n14481, n14482, n14484, n14485, n14486, n14487, n14488;
  wire n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496;
  wire n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504;
  wire n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512;
  wire n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520;
  wire n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528;
  wire n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14538;
  wire n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546;
  wire n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554;
  wire n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562;
  wire n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570;
  wire n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578;
  wire n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586;
  wire n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594;
  wire n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602;
  wire n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610;
  wire n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618;
  wire n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626;
  wire n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634;
  wire n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642;
  wire n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650;
  wire n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658;
  wire n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666;
  wire n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674;
  wire n14675, n14676, n14677, n14678, n14679, n14680, n14682, n14683;
  wire n14684, n14685, n14686, n14687, n14688, n14689, n14692, n14693;
  wire n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701;
  wire n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709;
  wire n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717;
  wire n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725;
  wire n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733;
  wire n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741;
  wire n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749;
  wire n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757;
  wire n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765;
  wire n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773;
  wire n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781;
  wire n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789;
  wire n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797;
  wire n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805;
  wire n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813;
  wire n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821;
  wire n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829;
  wire n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837;
  wire n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845;
  wire n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853;
  wire n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861;
  wire n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869;
  wire n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14878;
  wire n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886;
  wire n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894;
  wire n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902;
  wire n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910;
  wire n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918;
  wire n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928;
  wire n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936;
  wire n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944;
  wire n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952;
  wire n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960;
  wire n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968;
  wire n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976;
  wire n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984;
  wire n14985, n14986, n14989, n14990, n14991, n14992, n14993, n14994;
  wire n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002;
  wire n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010;
  wire n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018;
  wire n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026;
  wire n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034;
  wire n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042;
  wire n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050;
  wire n15051, n15052, n15053, n15054, n15055, n15057, n15058, n15059;
  wire n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067;
  wire n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075;
  wire n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083;
  wire n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091;
  wire n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099;
  wire n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107;
  wire n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115;
  wire n15116, n15117, n15118, n15119, n15122, n15123, n15124, n15125;
  wire n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133;
  wire n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141;
  wire n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149;
  wire n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157;
  wire n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165;
  wire n15166, n15167, n15168, n15169, n15172, n15173, n15174, n15175;
  wire n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183;
  wire n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191;
  wire n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199;
  wire n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207;
  wire n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215;
  wire n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223;
  wire n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231;
  wire n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15240;
  wire n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248;
  wire n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256;
  wire n15257, n15258, n15261, n15262, n15263, n15264, n15265, n15266;
  wire n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274;
  wire n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282;
  wire n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290;
  wire n15291, n15294, n15295, n15296, n15297, n15298, n15299, n15300;
  wire n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308;
  wire n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316;
  wire n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324;
  wire n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332;
  wire n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340;
  wire n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348;
  wire n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356;
  wire n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364;
  wire n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372;
  wire n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380;
  wire n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388;
  wire n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396;
  wire n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404;
  wire n15405, n15406, n15407, n15408, n15409, n15411, n15412, n15413;
  wire n15414, n15415, n15416, n15419, n15420, n15421, n15422, n15423;
  wire n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431;
  wire n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439;
  wire n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447;
  wire n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455;
  wire n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463;
  wire n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471;
  wire n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479;
  wire n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487;
  wire n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495;
  wire n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503;
  wire n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511;
  wire n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519;
  wire n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527;
  wire n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535;
  wire n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543;
  wire n15544, n15545, n15546, n15547, n15548, n15551, n15552, n15553;
  wire n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561;
  wire n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569;
  wire n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577;
  wire n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15586;
  wire n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594;
  wire n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602;
  wire n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610;
  wire n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618;
  wire n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626;
  wire n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634;
  wire n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642;
  wire n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650;
  wire n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658;
  wire n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666;
  wire n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674;
  wire n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682;
  wire n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690;
  wire n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698;
  wire n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706;
  wire n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714;
  wire n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722;
  wire n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730;
  wire n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738;
  wire n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746;
  wire n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754;
  wire n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763;
  wire n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771;
  wire n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779;
  wire n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787;
  wire n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795;
  wire n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803;
  wire n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811;
  wire n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819;
  wire n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827;
  wire n15828, n15829, n15830, n15831, n15834, n15835, n15836, n15837;
  wire n15838, n15839, n15840, n15841, n15842, n15843, n15846, n15847;
  wire n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855;
  wire n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863;
  wire n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871;
  wire n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879;
  wire n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887;
  wire n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895;
  wire n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903;
  wire n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911;
  wire n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919;
  wire n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928;
  wire n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936;
  wire n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944;
  wire n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952;
  wire n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960;
  wire n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968;
  wire n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976;
  wire n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984;
  wire n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992;
  wire n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000;
  wire n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008;
  wire n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016;
  wire n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024;
  wire n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032;
  wire n16033, n16034, n16035, n16036, n16037, n16040, n16041, n16042;
  wire n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050;
  wire n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058;
  wire n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066;
  wire n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074;
  wire n16075, n16077, n16078, n16079, n16080, n16081, n16082, n16083;
  wire n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091;
  wire n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099;
  wire n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107;
  wire n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115;
  wire n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123;
  wire n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131;
  wire n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139;
  wire n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147;
  wire n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155;
  wire n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163;
  wire n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171;
  wire n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179;
  wire n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187;
  wire n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195;
  wire n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203;
  wire n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211;
  wire n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219;
  wire n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16228;
  wire n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236;
  wire n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244;
  wire n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16254;
  wire n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262;
  wire n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270;
  wire n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278;
  wire n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286;
  wire n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294;
  wire n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302;
  wire n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310;
  wire n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318;
  wire n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326;
  wire n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334;
  wire n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342;
  wire n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350;
  wire n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358;
  wire n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366;
  wire n16367, n16368, n16370, n16371, n16372, n16373, n16374, n16375;
  wire n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383;
  wire n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391;
  wire n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399;
  wire n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407;
  wire n16408, n16409, n16410, n16411, n16414, n16415, n16416, n16417;
  wire n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425;
  wire n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433;
  wire n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441;
  wire n16442, n16443, n16444, n16445, n16446, n16447, n16450, n16451;
  wire n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459;
  wire n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467;
  wire n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475;
  wire n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483;
  wire n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491;
  wire n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499;
  wire n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507;
  wire n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515;
  wire n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524;
  wire n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532;
  wire n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540;
  wire n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548;
  wire n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556;
  wire n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564;
  wire n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572;
  wire n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580;
  wire n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588;
  wire n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596;
  wire n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604;
  wire n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612;
  wire n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620;
  wire n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628;
  wire n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636;
  wire n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644;
  wire n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652;
  wire n16653, n16654, n16655, n16656, n16657, n16659, n16660, n16661;
  wire n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669;
  wire n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677;
  wire n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685;
  wire n16686, n16687, n16688, n16691, n16692, n16693, n16694, n16695;
  wire n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703;
  wire n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711;
  wire n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719;
  wire n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727;
  wire n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735;
  wire n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743;
  wire n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751;
  wire n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759;
  wire n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767;
  wire n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775;
  wire n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783;
  wire n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791;
  wire n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800;
  wire n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808;
  wire n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816;
  wire n16817, n16820, n16821, n16822, n16823, n16824, n16825, n16826;
  wire n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834;
  wire n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842;
  wire n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850;
  wire n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858;
  wire n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866;
  wire n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874;
  wire n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882;
  wire n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890;
  wire n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898;
  wire n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906;
  wire n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914;
  wire n16915, n16916, n16918, n16919, n16920, n16921, n16922, n16923;
  wire n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931;
  wire n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939;
  wire n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947;
  wire n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955;
  wire n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963;
  wire n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971;
  wire n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979;
  wire n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987;
  wire n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995;
  wire n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003;
  wire n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011;
  wire n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019;
  wire n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027;
  wire n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035;
  wire n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043;
  wire n17044, n17045, n17046, n17048, n17049, n17050, n17051, n17052;
  wire n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060;
  wire n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068;
  wire n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076;
  wire n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084;
  wire n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092;
  wire n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100;
  wire n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108;
  wire n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116;
  wire n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124;
  wire n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132;
  wire n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140;
  wire n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148;
  wire n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156;
  wire n17157, n17158, n17160, n17161, n17162, n17163, n17164, n17165;
  wire n17166, n17169, n17170, n17171, n17172, n17173, n17174, n17175;
  wire n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183;
  wire n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191;
  wire n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199;
  wire n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207;
  wire n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215;
  wire n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223;
  wire n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231;
  wire n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239;
  wire n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247;
  wire n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255;
  wire n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263;
  wire n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271;
  wire n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17280;
  wire n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288;
  wire n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296;
  wire n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304;
  wire n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312;
  wire n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320;
  wire n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328;
  wire n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336;
  wire n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344;
  wire n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352;
  wire n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360;
  wire n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368;
  wire n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376;
  wire n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384;
  wire n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392;
  wire n17393, n17394, n17396, n17397, n17398, n17399, n17400, n17401;
  wire n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411;
  wire n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419;
  wire n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427;
  wire n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435;
  wire n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443;
  wire n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451;
  wire n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459;
  wire n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467;
  wire n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475;
  wire n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483;
  wire n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491;
  wire n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499;
  wire n17500, n17501, n17503, n17504, n17505, n17506, n17507, n17508;
  wire n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516;
  wire n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524;
  wire n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532;
  wire n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540;
  wire n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548;
  wire n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556;
  wire n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564;
  wire n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572;
  wire n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580;
  wire n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588;
  wire n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596;
  wire n17597, n17598, n17599, n17600, n17601, n17603, n17604, n17605;
  wire n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613;
  wire n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621;
  wire n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629;
  wire n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637;
  wire n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645;
  wire n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653;
  wire n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661;
  wire n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669;
  wire n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677;
  wire n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685;
  wire n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693;
  wire n17694, n17695, n17696, n17697, n17698, n17699, n17701, n17702;
  wire n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710;
  wire n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718;
  wire n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726;
  wire n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734;
  wire n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742;
  wire n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750;
  wire n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758;
  wire n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766;
  wire n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774;
  wire n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782;
  wire n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790;
  wire n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799;
  wire n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807;
  wire n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815;
  wire n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823;
  wire n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831;
  wire n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839;
  wire n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847;
  wire n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855;
  wire n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863;
  wire n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871;
  wire n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879;
  wire n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888;
  wire n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896;
  wire n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904;
  wire n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912;
  wire n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920;
  wire n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928;
  wire n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936;
  wire n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944;
  wire n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952;
  wire n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960;
  wire n17961, n17962, n17963, n17964, n17965, n17967, n17968, n17969;
  wire n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977;
  wire n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985;
  wire n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993;
  wire n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001;
  wire n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009;
  wire n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017;
  wire n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025;
  wire n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033;
  wire n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041;
  wire n18042, n18043, n18044, n18046, n18047, n18048, n18049, n18050;
  wire n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058;
  wire n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066;
  wire n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074;
  wire n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082;
  wire n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090;
  wire n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098;
  wire n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106;
  wire n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114;
  wire n18115, n18116, n18117, n18118, n18119, n18120, n18122, n18123;
  wire n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131;
  wire n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139;
  wire n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147;
  wire n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155;
  wire n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163;
  wire n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171;
  wire n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179;
  wire n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187;
  wire n18188, n18189, n18190, n18191, n18193, n18194, n18195, n18196;
  wire n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204;
  wire n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212;
  wire n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220;
  wire n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228;
  wire n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236;
  wire n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244;
  wire n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252;
  wire n18253, n18254, n18256, n18257, n18258, n18259, n18260, n18261;
  wire n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269;
  wire n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277;
  wire n18278, n18279, n18280, n18283, n18284, n18285, n18286, n18287;
  wire n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295;
  wire n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303;
  wire n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311;
  wire n18312, n18314, n18315, n18316, n18317, n18318, n18319, n18320;
  wire n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328;
  wire n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336;
  wire n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344;
  wire n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352;
  wire n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360;
  wire n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368;
  wire n18369, n18371, n18372, n18373, n18374, n18375, n18376, n18377;
  wire n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385;
  wire n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393;
  wire n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401;
  wire n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409;
  wire n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417;
  wire n18418, n18419, n18421, n18422, n18423, n18424, n18425, n18426;
  wire n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434;
  wire n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442;
  wire n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450;
  wire n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458;
  wire n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466;
  wire n18467, n18469, n18470, n18471, n18472, n18473, n18474, n18475;
  wire n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483;
  wire n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491;
  wire n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499;
  wire n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507;
  wire n18508, n18509, n18510, n18511, n18513, n18514, n18515, n18516;
  wire n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524;
  wire n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532;
  wire n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540;
  wire n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18549;
  wire n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557;
  wire n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565;
  wire n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573;
  wire n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581;
  wire n18582, n18584, n18585, n18586, n18587, n18588, n18589, n18590;
  wire n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598;
  wire n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606;
  wire n18607, n18608, n18609, n18610, n18611, n18613, n18614, n18615;
  wire n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623;
  wire n18624, n18625, n18626, n18627, n18628, n18629, n18631, n18632;
  wire n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640;
  wire n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648;
  wire n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657;
  wire n18658, n18659, n18661, n18662, n18663, n18664, n18665, n18666;
  wire n18667, n18668, n18670, n18671, n18672, n18673, n18674, n18676;
  wire n_4, n_6, n_7, n_8, n_9, n_11, n_12, n_13;
  wire n_14, n_15, n_17, n_18, n_19, n_20, n_21, n_22;
  wire n_23, n_24, n_25, n_26, n_27, n_29, n_30, n_31;
  wire n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_256, n_257, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555;
  wire n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595;
  wire n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603;
  wire n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611;
  wire n_612, n_613, n_614, n_615, n_616, n_617, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644;
  wire n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
  wire n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724;
  wire n_725, n_726, n_727, n_728, n_730, n_731, n_732, n_733;
  wire n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757;
  wire n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765;
  wire n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781;
  wire n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789;
  wire n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813;
  wire n_814, n_816, n_817, n_818, n_819, n_820, n_821, n_822;
  wire n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830;
  wire n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838;
  wire n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846;
  wire n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
  wire n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870;
  wire n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878;
  wire n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902;
  wire n_903, n_904, n_905, n_906, n_907, n_908, n_910, n_911;
  wire n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919;
  wire n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927;
  wire n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935;
  wire n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943;
  wire n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_963, n_964, n_965, n_966, n_967, n_968;
  wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
  wire n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984;
  wire n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016;
  wire n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048;
  wire n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056;
  wire n_1057, n_1058, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065;
  wire n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073;
  wire n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089;
  wire n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097;
  wire n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105;
  wire n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113;
  wire n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121;
  wire n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129;
  wire n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137;
  wire n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1152, n_1153, n_1154;
  wire n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186;
  wire n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202;
  wire n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210;
  wire n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218;
  wire n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226;
  wire n_1227, n_1228, n_1229, n_1231, n_1232, n_1233, n_1234, n_1235;
  wire n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243;
  wire n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267;
  wire n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275;
  wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
  wire n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307;
  wire n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315;
  wire n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323;
  wire n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
  wire n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347;
  wire n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355;
  wire n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1388, n_1389, n_1390, n_1392, n_1393, n_1394, n_1395, n_1396;
  wire n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404;
  wire n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412;
  wire n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420;
  wire n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428;
  wire n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436;
  wire n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444;
  wire n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452;
  wire n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460;
  wire n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468;
  wire n_1469, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477;
  wire n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485;
  wire n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501;
  wire n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509;
  wire n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
  wire n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565;
  wire n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573;
  wire n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581;
  wire n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589;
  wire n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597;
  wire n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605;
  wire n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1627, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638;
  wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654;
  wire n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662;
  wire n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670;
  wire n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678;
  wire n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711;
  wire n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719;
  wire n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727;
  wire n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
  wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872;
  wire n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880;
  wire n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888;
  wire n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896;
  wire n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920;
  wire n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928;
  wire n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936;
  wire n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1958, n_1959, n_1960, n_1961;
  wire n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969;
  wire n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977;
  wire n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985;
  wire n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993;
  wire n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001;
  wire n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009;
  wire n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017;
  wire n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025;
  wire n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057;
  wire n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073;
  wire n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081;
  wire n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098;
  wire n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106;
  wire n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114;
  wire n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122;
  wire n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130;
  wire n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138;
  wire n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146;
  wire n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154;
  wire n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162;
  wire n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170;
  wire n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186;
  wire n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194;
  wire n_2195, n_2196, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203;
  wire n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211;
  wire n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219;
  wire n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227;
  wire n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235;
  wire n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243;
  wire n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251;
  wire n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259;
  wire n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267;
  wire n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275;
  wire n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283;
  wire n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291;
  wire n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299;
  wire n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307;
  wire n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315;
  wire n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323;
  wire n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331;
  wire n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339;
  wire n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347;
  wire n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355;
  wire n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363;
  wire n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371;
  wire n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379;
  wire n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387;
  wire n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395;
  wire n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403;
  wire n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411;
  wire n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419;
  wire n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2435, n_2436;
  wire n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468;
  wire n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476;
  wire n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484;
  wire n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492;
  wire n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500;
  wire n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508;
  wire n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516;
  wire n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524;
  wire n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2532, n_2533;
  wire n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541;
  wire n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549;
  wire n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557;
  wire n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565;
  wire n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573;
  wire n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581;
  wire n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589;
  wire n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597;
  wire n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605;
  wire n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613;
  wire n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621;
  wire n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629;
  wire n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637;
  wire n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645;
  wire n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653;
  wire n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661;
  wire n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669;
  wire n_2670, n_2671, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678;
  wire n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686;
  wire n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694;
  wire n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702;
  wire n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710;
  wire n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718;
  wire n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726;
  wire n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734;
  wire n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742;
  wire n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750;
  wire n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758;
  wire n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782;
  wire n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790;
  wire n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798;
  wire n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806;
  wire n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814;
  wire n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822;
  wire n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830;
  wire n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838;
  wire n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847;
  wire n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855;
  wire n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863;
  wire n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871;
  wire n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879;
  wire n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887;
  wire n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895;
  wire n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903;
  wire n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911;
  wire n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919;
  wire n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927;
  wire n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935;
  wire n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943;
  wire n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951;
  wire n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959;
  wire n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967;
  wire n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975;
  wire n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983;
  wire n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991;
  wire n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999;
  wire n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007;
  wire n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015;
  wire n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023;
  wire n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031;
  wire n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039;
  wire n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048;
  wire n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056;
  wire n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064;
  wire n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072;
  wire n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080;
  wire n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3089;
  wire n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097;
  wire n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105;
  wire n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113;
  wire n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121;
  wire n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129;
  wire n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137;
  wire n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145;
  wire n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153;
  wire n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161;
  wire n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169;
  wire n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177;
  wire n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185;
  wire n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193;
  wire n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201;
  wire n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209;
  wire n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217;
  wire n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225;
  wire n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233;
  wire n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241;
  wire n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249;
  wire n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257;
  wire n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265;
  wire n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273;
  wire n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281;
  wire n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289;
  wire n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297;
  wire n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306;
  wire n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314;
  wire n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322;
  wire n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330;
  wire n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338;
  wire n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346;
  wire n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354;
  wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362;
  wire n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370;
  wire n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378;
  wire n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386;
  wire n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394;
  wire n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402;
  wire n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410;
  wire n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418;
  wire n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426;
  wire n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434;
  wire n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442;
  wire n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450;
  wire n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458;
  wire n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, n_3466;
  wire n_3467, n_3468, n_3469, n_3470, n_3471, n_3473, n_3474, n_3475;
  wire n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483;
  wire n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491;
  wire n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499;
  wire n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507;
  wire n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515;
  wire n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523;
  wire n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531;
  wire n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539;
  wire n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547;
  wire n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555;
  wire n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563;
  wire n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571;
  wire n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579;
  wire n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587;
  wire n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595;
  wire n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603;
  wire n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611;
  wire n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619;
  wire n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627;
  wire n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635;
  wire n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643;
  wire n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651;
  wire n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659;
  wire n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667;
  wire n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675;
  wire n_3676, n_3677, n_3678, n_3679, n_3681, n_3682, n_3683, n_3684;
  wire n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692;
  wire n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700;
  wire n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708;
  wire n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716;
  wire n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724;
  wire n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732;
  wire n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, n_3740;
  wire n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748;
  wire n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756;
  wire n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764;
  wire n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772;
  wire n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780;
  wire n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788;
  wire n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796;
  wire n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804;
  wire n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3813;
  wire n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821;
  wire n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829;
  wire n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837;
  wire n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845;
  wire n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, n_3853;
  wire n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861;
  wire n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869;
  wire n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877;
  wire n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885;
  wire n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893;
  wire n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901;
  wire n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909;
  wire n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917;
  wire n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, n_3925;
  wire n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, n_3933;
  wire n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941;
  wire n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949;
  wire n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957;
  wire n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965;
  wire n_3966, n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973;
  wire n_3974, n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981;
  wire n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989;
  wire n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997;
  wire n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005;
  wire n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013;
  wire n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021;
  wire n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029;
  wire n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037;
  wire n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045;
  wire n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053;
  wire n_4054, n_4055, n_4056, n_4058, n_4059, n_4060, n_4061, n_4062;
  wire n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070;
  wire n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078;
  wire n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086;
  wire n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094;
  wire n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102;
  wire n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110;
  wire n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118;
  wire n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126;
  wire n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134;
  wire n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142;
  wire n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150;
  wire n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158;
  wire n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166;
  wire n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174;
  wire n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182;
  wire n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190;
  wire n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198;
  wire n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206;
  wire n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214;
  wire n_4215, n_4216, n_4217, n_4219, n_4220, n_4221, n_4222, n_4223;
  wire n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231;
  wire n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239;
  wire n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247;
  wire n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255;
  wire n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263;
  wire n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271;
  wire n_4272, n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279;
  wire n_4280, n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287;
  wire n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295;
  wire n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303;
  wire n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311;
  wire n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319;
  wire n_4320, n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327;
  wire n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335;
  wire n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343;
  wire n_4344, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351;
  wire n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359;
  wire n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367;
  wire n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375;
  wire n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383;
  wire n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391;
  wire n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399;
  wire n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407;
  wire n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416;
  wire n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424;
  wire n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432;
  wire n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440;
  wire n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448;
  wire n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456;
  wire n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464;
  wire n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472;
  wire n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480;
  wire n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488;
  wire n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496;
  wire n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504;
  wire n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512;
  wire n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520;
  wire n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528;
  wire n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536;
  wire n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544;
  wire n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552;
  wire n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560;
  wire n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568;
  wire n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576;
  wire n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584;
  wire n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592;
  wire n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600;
  wire n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608;
  wire n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616;
  wire n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4625;
  wire n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633;
  wire n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641;
  wire n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649;
  wire n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657;
  wire n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665;
  wire n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673;
  wire n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681;
  wire n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689;
  wire n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697;
  wire n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705;
  wire n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713;
  wire n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721;
  wire n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728, n_4729;
  wire n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737;
  wire n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745;
  wire n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752, n_4753;
  wire n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760, n_4761;
  wire n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768, n_4769;
  wire n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777;
  wire n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785;
  wire n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4793;
  wire n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800, n_4801;
  wire n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809;
  wire n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817;
  wire n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825;
  wire n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832, n_4833;
  wire n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840, n_4841;
  wire n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848, n_4849;
  wire n_4850, n_4851, n_4852, n_4853, n_4854, n_4856, n_4857, n_4858;
  wire n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866;
  wire n_4867, n_4868, n_4869, n_4870, n_4871, n_4872, n_4873, n_4874;
  wire n_4875, n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882;
  wire n_4883, n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4890;
  wire n_4891, n_4892, n_4893, n_4894, n_4895, n_4896, n_4897, n_4898;
  wire n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906;
  wire n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914;
  wire n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922;
  wire n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930;
  wire n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938;
  wire n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946;
  wire n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954;
  wire n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962;
  wire n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970;
  wire n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978;
  wire n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986;
  wire n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994;
  wire n_4995, n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002;
  wire n_5003, n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010;
  wire n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018;
  wire n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026;
  wire n_5027, n_5028, n_5029, n_5030, n_5032, n_5033, n_5034, n_5035;
  wire n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043;
  wire n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051;
  wire n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059;
  wire n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067;
  wire n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075;
  wire n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083;
  wire n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091;
  wire n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099;
  wire n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107;
  wire n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115;
  wire n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123;
  wire n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131;
  wire n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139;
  wire n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147;
  wire n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155;
  wire n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163;
  wire n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171;
  wire n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179;
  wire n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187;
  wire n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195;
  wire n_5196, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204;
  wire n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, n_5212;
  wire n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220;
  wire n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228;
  wire n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236;
  wire n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244;
  wire n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252;
  wire n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260;
  wire n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268;
  wire n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276;
  wire n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283, n_5284;
  wire n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291, n_5292;
  wire n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299, n_5300;
  wire n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307, n_5308;
  wire n_5309, n_5310, n_5311, n_5312, n_5313, n_5314, n_5315, n_5316;
  wire n_5317, n_5318, n_5319, n_5320, n_5321, n_5322, n_5323, n_5324;
  wire n_5325, n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5332;
  wire n_5333, n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5340;
  wire n_5341, n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348;
  wire n_5349, n_5350, n_5351, n_5352, n_5353, n_5354, n_5355, n_5356;
  wire n_5357, n_5358, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364;
  wire n_5365, n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372;
  wire n_5373, n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380;
  wire n_5381, n_5382, n_5383, n_5384, n_5385, n_5387, n_5388, n_5389;
  wire n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397;
  wire n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405;
  wire n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413;
  wire n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421;
  wire n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429;
  wire n_5430, n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, n_5437;
  wire n_5438, n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445;
  wire n_5446, n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453;
  wire n_5454, n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461;
  wire n_5462, n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469;
  wire n_5470, n_5471, n_5472, n_5473, n_5474, n_5475, n_5476, n_5477;
  wire n_5478, n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485;
  wire n_5486, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493;
  wire n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501;
  wire n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509;
  wire n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517;
  wire n_5518, n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525;
  wire n_5526, n_5527, n_5528, n_5529, n_5530, n_5531, n_5532, n_5533;
  wire n_5534, n_5535, n_5536, n_5537, n_5538, n_5539, n_5540, n_5541;
  wire n_5542, n_5543, n_5544, n_5545, n_5546, n_5547, n_5548, n_5549;
  wire n_5550, n_5551, n_5552, n_5553, n_5554, n_5555, n_5556, n_5557;
  wire n_5558, n_5559, n_5560, n_5561, n_5562, n_5563, n_5564, n_5565;
  wire n_5566, n_5567, n_5568, n_5569, n_5570, n_5571, n_5572, n_5573;
  wire n_5574, n_5575, n_5576, n_5577, n_5578, n_5579, n_5580, n_5581;
  wire n_5582, n_5583, n_5584, n_5585, n_5586, n_5587, n_5588, n_5589;
  wire n_5590, n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597;
  wire n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605;
  wire n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613;
  wire n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621;
  wire n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629;
  wire n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637;
  wire n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645;
  wire n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653;
  wire n_5654, n_5655, n_5656, n_5657, n_5659, n_5660, n_5661, n_5662;
  wire n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669, n_5670;
  wire n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677, n_5678;
  wire n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686;
  wire n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5694;
  wire n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702;
  wire n_5703, n_5704, n_5705, n_5706, n_5707, n_5708, n_5709, n_5710;
  wire n_5711, n_5712, n_5713, n_5714, n_5715, n_5716, n_5717, n_5718;
  wire n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726;
  wire n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734;
  wire n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742;
  wire n_5743, n_5744, n_5745, n_5746, n_5747, n_5748, n_5749, n_5750;
  wire n_5751, n_5752, n_5753, n_5754, n_5755, n_5756, n_5757, n_5758;
  wire n_5759, n_5760, n_5761, n_5762, n_5763, n_5764, n_5765, n_5766;
  wire n_5767, n_5768, n_5769, n_5770, n_5771, n_5772, n_5773, n_5774;
  wire n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781, n_5782;
  wire n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789, n_5790;
  wire n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797, n_5798;
  wire n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806;
  wire n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813, n_5814;
  wire n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822;
  wire n_5823, n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830;
  wire n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838;
  wire n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846;
  wire n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854;
  wire n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861, n_5862;
  wire n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869, n_5870;
  wire n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877, n_5878;
  wire n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885, n_5886;
  wire n_5887, n_5888, n_5889, n_5890, n_5891, n_5893, n_5894, n_5895;
  wire n_5896, n_5897, n_5898, n_5899, n_5900, n_5901, n_5902, n_5903;
  wire n_5904, n_5905, n_5906, n_5907, n_5908, n_5909, n_5910, n_5911;
  wire n_5912, n_5913, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919;
  wire n_5920, n_5921, n_5922, n_5923, n_5924, n_5925, n_5926, n_5927;
  wire n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935;
  wire n_5936, n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943;
  wire n_5944, n_5945, n_5946, n_5947, n_5948, n_5949, n_5950, n_5951;
  wire n_5952, n_5953, n_5954, n_5955, n_5956, n_5957, n_5958, n_5959;
  wire n_5960, n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967;
  wire n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975;
  wire n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983;
  wire n_5984, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991;
  wire n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999;
  wire n_6000, n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007;
  wire n_6008, n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015;
  wire n_6016, n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023;
  wire n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031;
  wire n_6032, n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039;
  wire n_6040, n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047;
  wire n_6048, n_6049, n_6050, n_6051, n_6052, n_6054, n_6055, n_6056;
  wire n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064;
  wire n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072;
  wire n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080;
  wire n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087, n_6088;
  wire n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095, n_6096;
  wire n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104;
  wire n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112;
  wire n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120;
  wire n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128;
  wire n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136;
  wire n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144;
  wire n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152;
  wire n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160;
  wire n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168;
  wire n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176;
  wire n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184;
  wire n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192;
  wire n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200;
  wire n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208;
  wire n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216;
  wire n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224;
  wire n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232;
  wire n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240;
  wire n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247, n_6248;
  wire n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256;
  wire n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263, n_6264;
  wire n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271, n_6272;
  wire n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279, n_6280;
  wire n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287, n_6288;
  wire n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295, n_6296;
  wire n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303, n_6304;
  wire n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311, n_6312;
  wire n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319, n_6320;
  wire n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328;
  wire n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336;
  wire n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344;
  wire n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6352;
  wire n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359, n_6360;
  wire n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367, n_6368;
  wire n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376;
  wire n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384;
  wire n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392;
  wire n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400;
  wire n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408;
  wire n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416;
  wire n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424;
  wire n_6425, n_6426, n_6427, n_6428, n_6429, n_6430, n_6431, n_6432;
  wire n_6433, n_6434, n_6435, n_6436, n_6437, n_6438, n_6439, n_6440;
  wire n_6442, n_6443, n_6444, n_6445, n_6446, n_6447, n_6448, n_6449;
  wire n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457;
  wire n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, n_6465;
  wire n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472, n_6473;
  wire n_6474, n_6475, n_6476, n_6477, n_6478, n_6479, n_6480, n_6481;
  wire n_6482, n_6483, n_6484, n_6485, n_6486, n_6487, n_6488, n_6489;
  wire n_6490, n_6491, n_6492, n_6493, n_6494, n_6495, n_6496, n_6497;
  wire n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504, n_6505;
  wire n_6506, n_6507, n_6508, n_6509, n_6510, n_6511, n_6512, n_6513;
  wire n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520, n_6521;
  wire n_6522, n_6523, n_6524, n_6525, n_6526, n_6527, n_6528, n_6529;
  wire n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536, n_6537;
  wire n_6538, n_6539, n_6540, n_6541, n_6542, n_6543, n_6544, n_6545;
  wire n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6552, n_6553;
  wire n_6554, n_6555, n_6556, n_6557, n_6558, n_6559, n_6560, n_6561;
  wire n_6562, n_6563, n_6564, n_6565, n_6566, n_6567, n_6568, n_6569;
  wire n_6570, n_6571, n_6572, n_6573, n_6574, n_6575, n_6576, n_6577;
  wire n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6585;
  wire n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592, n_6593;
  wire n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601;
  wire n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6609, n_6610;
  wire n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617, n_6618;
  wire n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6625, n_6626;
  wire n_6627, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6634;
  wire n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641, n_6642;
  wire n_6643, n_6644, n_6645, n_6646, n_6647, n_6648, n_6649, n_6650;
  wire n_6651, n_6652, n_6653, n_6654, n_6655, n_6656, n_6657, n_6658;
  wire n_6659, n_6660, n_6661, n_6662, n_6663, n_6664, n_6665, n_6666;
  wire n_6667, n_6668, n_6669, n_6670, n_6671, n_6672, n_6673, n_6674;
  wire n_6675, n_6676, n_6677, n_6678, n_6679, n_6680, n_6681, n_6682;
  wire n_6683, n_6684, n_6685, n_6686, n_6687, n_6688, n_6689, n_6690;
  wire n_6691, n_6692, n_6693, n_6694, n_6695, n_6696, n_6697, n_6698;
  wire n_6699, n_6700, n_6701, n_6702, n_6703, n_6704, n_6705, n_6706;
  wire n_6707, n_6708, n_6709, n_6710, n_6711, n_6712, n_6713, n_6714;
  wire n_6715, n_6716, n_6717, n_6718, n_6719, n_6720, n_6721, n_6722;
  wire n_6723, n_6724, n_6725, n_6726, n_6727, n_6728, n_6729, n_6730;
  wire n_6731, n_6732, n_6733, n_6734, n_6735, n_6736, n_6737, n_6738;
  wire n_6739, n_6740, n_6741, n_6742, n_6743, n_6744, n_6745, n_6746;
  wire n_6747, n_6748, n_6749, n_6750, n_6751, n_6752, n_6753, n_6754;
  wire n_6755, n_6756, n_6757, n_6758, n_6759, n_6760, n_6761, n_6762;
  wire n_6763, n_6764, n_6765, n_6766, n_6767, n_6768, n_6769, n_6770;
  wire n_6771, n_6772, n_6773, n_6774, n_6775, n_6776, n_6777, n_6778;
  wire n_6779, n_6780, n_6781, n_6782, n_6783, n_6784, n_6785, n_6786;
  wire n_6787, n_6788, n_6789, n_6790, n_6791, n_6792, n_6793, n_6794;
  wire n_6795, n_6796, n_6797, n_6798, n_6799, n_6800, n_6801, n_6802;
  wire n_6803, n_6804, n_6805, n_6806, n_6807, n_6808, n_6809, n_6810;
  wire n_6811, n_6812, n_6813, n_6814, n_6815, n_6816, n_6817, n_6818;
  wire n_6819, n_6820, n_6821, n_6822, n_6823, n_6824, n_6825, n_6826;
  wire n_6827, n_6828, n_6829, n_6830, n_6831, n_6832, n_6833, n_6834;
  wire n_6835, n_6836, n_6837, n_6838, n_6839, n_6840, n_6841, n_6842;
  wire n_6843, n_6844, n_6845, n_6846, n_6847, n_6848, n_6849, n_6850;
  wire n_6851, n_6852, n_6853, n_6854, n_6855, n_6856, n_6857, n_6858;
  wire n_6859, n_6860, n_6861, n_6862, n_6863, n_6864, n_6865, n_6866;
  wire n_6867, n_6868, n_6869, n_6870, n_6871, n_6872, n_6873, n_6874;
  wire n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881, n_6882;
  wire n_6883, n_6884, n_6885, n_6886, n_6887, n_6888, n_6889, n_6890;
  wire n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6898;
  wire n_6899, n_6900, n_6901, n_6902, n_6903, n_6904, n_6905, n_6906;
  wire n_6907, n_6908, n_6909, n_6910, n_6911, n_6912, n_6913, n_6914;
  wire n_6915, n_6916, n_6917, n_6918, n_6919, n_6920, n_6921, n_6922;
  wire n_6923, n_6924, n_6925, n_6926, n_6927, n_6928, n_6929, n_6930;
  wire n_6931, n_6932, n_6933, n_6934, n_6935, n_6936, n_6937, n_6938;
  wire n_6939, n_6940, n_6941, n_6942, n_6943, n_6944, n_6945, n_6946;
  wire n_6947, n_6948, n_6949, n_6950, n_6951, n_6952, n_6953, n_6954;
  wire n_6955, n_6956, n_6957, n_6958, n_6959, n_6961, n_6962, n_6963;
  wire n_6964, n_6965, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971;
  wire n_6972, n_6973, n_6974, n_6975, n_6976, n_6977, n_6978, n_6979;
  wire n_6980, n_6981, n_6982, n_6983, n_6984, n_6985, n_6986, n_6987;
  wire n_6988, n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995;
  wire n_6996, n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, n_7003;
  wire n_7004, n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011;
  wire n_7012, n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019;
  wire n_7020, n_7021, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027;
  wire n_7028, n_7029, n_7030, n_7031, n_7032, n_7033, n_7034, n_7035;
  wire n_7036, n_7037, n_7038, n_7039, n_7040, n_7041, n_7042, n_7043;
  wire n_7044, n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7051;
  wire n_7052, n_7053, n_7054, n_7055, n_7056, n_7057, n_7058, n_7059;
  wire n_7060, n_7061, n_7062, n_7063, n_7064, n_7065, n_7066, n_7067;
  wire n_7068, n_7069, n_7070, n_7071, n_7072, n_7073, n_7074, n_7075;
  wire n_7076, n_7077, n_7078, n_7079, n_7080, n_7081, n_7082, n_7083;
  wire n_7084, n_7085, n_7086, n_7087, n_7088, n_7089, n_7090, n_7091;
  wire n_7092, n_7093, n_7095, n_7096, n_7097, n_7098, n_7099, n_7100;
  wire n_7101, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108;
  wire n_7109, n_7110, n_7111, n_7112, n_7113, n_7114, n_7115, n_7116;
  wire n_7117, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123, n_7124;
  wire n_7125, n_7126, n_7127, n_7128, n_7129, n_7130, n_7131, n_7132;
  wire n_7133, n_7134, n_7135, n_7136, n_7137, n_7138, n_7139, n_7140;
  wire n_7141, n_7142, n_7143, n_7144, n_7145, n_7146, n_7147, n_7148;
  wire n_7149, n_7150, n_7151, n_7152, n_7153, n_7154, n_7155, n_7156;
  wire n_7157, n_7158, n_7159, n_7160, n_7161, n_7162, n_7163, n_7164;
  wire n_7165, n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172;
  wire n_7173, n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180;
  wire n_7181, n_7182, n_7183, n_7184, n_7185, n_7186, n_7187, n_7188;
  wire n_7189, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195, n_7196;
  wire n_7197, n_7198, n_7199, n_7200, n_7201, n_7202, n_7203, n_7204;
  wire n_7205, n_7206, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212;
  wire n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220;
  wire n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228;
  wire n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236;
  wire n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7243, n_7244;
  wire n_7245, n_7246, n_7247, n_7248, n_7249, n_7250, n_7251, n_7252;
  wire n_7253, n_7254, n_7255, n_7256, n_7257, n_7258, n_7259, n_7260;
  wire n_7261, n_7262, n_7263, n_7264, n_7265, n_7266, n_7267, n_7268;
  wire n_7269, n_7270, n_7271, n_7272, n_7273, n_7274, n_7275, n_7276;
  wire n_7277, n_7278, n_7279, n_7280, n_7281, n_7282, n_7283, n_7284;
  wire n_7285, n_7286, n_7287, n_7288, n_7289, n_7290, n_7291, n_7292;
  wire n_7293, n_7294, n_7295, n_7296, n_7297, n_7298, n_7299, n_7300;
  wire n_7301, n_7302, n_7303, n_7304, n_7305, n_7306, n_7307, n_7308;
  wire n_7309, n_7310, n_7311, n_7312, n_7313, n_7314, n_7315, n_7316;
  wire n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7323, n_7324;
  wire n_7325, n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332;
  wire n_7333, n_7334, n_7335, n_7336, n_7337, n_7338, n_7339, n_7340;
  wire n_7341, n_7342, n_7343, n_7344, n_7345, n_7346, n_7347, n_7348;
  wire n_7349, n_7350, n_7351, n_7352, n_7353, n_7354, n_7355, n_7356;
  wire n_7357, n_7358, n_7359, n_7360, n_7361, n_7362, n_7363, n_7364;
  wire n_7365, n_7366, n_7367, n_7368, n_7369, n_7370, n_7371, n_7372;
  wire n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, n_7380;
  wire n_7381, n_7382, n_7383, n_7384, n_7385, n_7386, n_7387, n_7388;
  wire n_7389, n_7390, n_7391, n_7392, n_7393, n_7394, n_7395, n_7396;
  wire n_7397, n_7398, n_7399, n_7400, n_7401, n_7402, n_7403, n_7404;
  wire n_7405, n_7406, n_7407, n_7408, n_7409, n_7410, n_7412, n_7413;
  wire n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7421;
  wire n_7422, n_7423, n_7424, n_7425, n_7426, n_7427, n_7428, n_7429;
  wire n_7430, n_7431, n_7432, n_7433, n_7434, n_7435, n_7436, n_7437;
  wire n_7438, n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445;
  wire n_7446, n_7447, n_7448, n_7449, n_7450, n_7451, n_7452, n_7453;
  wire n_7454, n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461;
  wire n_7462, n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469;
  wire n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477;
  wire n_7478, n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485;
  wire n_7486, n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493;
  wire n_7494, n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501;
  wire n_7502, n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509;
  wire n_7510, n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517;
  wire n_7518, n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525;
  wire n_7526, n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533;
  wire n_7534, n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541;
  wire n_7542, n_7543, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549;
  wire n_7550, n_7551, n_7552, n_7553, n_7554, n_7555, n_7556, n_7557;
  wire n_7558, n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565;
  wire n_7566, n_7567, n_7568, n_7569, n_7570, n_7571, n_7572, n_7573;
  wire n_7574, n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581;
  wire n_7582, n_7583, n_7584, n_7585, n_7586, n_7587, n_7588, n_7589;
  wire n_7590, n_7591, n_7592, n_7593, n_7594, n_7595, n_7596, n_7597;
  wire n_7598, n_7599, n_7600, n_7601, n_7602, n_7603, n_7604, n_7605;
  wire n_7606, n_7607, n_7608, n_7609, n_7610, n_7611, n_7612, n_7613;
  wire n_7614, n_7615, n_7617, n_7618, n_7619, n_7620, n_7621, n_7622;
  wire n_7623, n_7624, n_7625, n_7626, n_7627, n_7628, n_7629, n_7630;
  wire n_7631, n_7632, n_7633, n_7634, n_7635, n_7636, n_7637, n_7638;
  wire n_7639, n_7640, n_7641, n_7642, n_7643, n_7644, n_7645, n_7646;
  wire n_7647, n_7648, n_7649, n_7650, n_7651, n_7652, n_7653, n_7654;
  wire n_7655, n_7656, n_7657, n_7658, n_7659, n_7660, n_7661, n_7662;
  wire n_7663, n_7664, n_7665, n_7666, n_7667, n_7668, n_7669, n_7670;
  wire n_7671, n_7672, n_7673, n_7674, n_7675, n_7676, n_7677, n_7678;
  wire n_7679, n_7680, n_7681, n_7682, n_7683, n_7684, n_7685, n_7686;
  wire n_7687, n_7688, n_7689, n_7690, n_7691, n_7692, n_7693, n_7694;
  wire n_7695, n_7696, n_7697, n_7698, n_7699, n_7700, n_7701, n_7702;
  wire n_7703, n_7704, n_7705, n_7706, n_7707, n_7708, n_7709, n_7710;
  wire n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717, n_7718;
  wire n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726;
  wire n_7727, n_7728, n_7729, n_7730, n_7731, n_7732, n_7733, n_7734;
  wire n_7735, n_7736, n_7737, n_7738, n_7739, n_7740, n_7741, n_7742;
  wire n_7743, n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750;
  wire n_7751, n_7752, n_7753, n_7754, n_7755, n_7756, n_7757, n_7758;
  wire n_7759, n_7760, n_7761, n_7762, n_7763, n_7764, n_7765, n_7766;
  wire n_7767, n_7768, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774;
  wire n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781, n_7782;
  wire n_7783, n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790;
  wire n_7791, n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798;
  wire n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7806;
  wire n_7807, n_7808, n_7809, n_7810, n_7811, n_7812, n_7813, n_7814;
  wire n_7815, n_7816, n_7817, n_7818, n_7819, n_7820, n_7821, n_7822;
  wire n_7823, n_7824, n_7825, n_7826, n_7827, n_7828, n_7829, n_7830;
  wire n_7831, n_7832, n_7833, n_7834, n_7835, n_7836, n_7837, n_7838;
  wire n_7839, n_7840, n_7841, n_7842, n_7843, n_7844, n_7845, n_7846;
  wire n_7847, n_7848, n_7849, n_7850, n_7851, n_7852, n_7853, n_7854;
  wire n_7855, n_7856, n_7857, n_7858, n_7859, n_7860, n_7861, n_7862;
  wire n_7863, n_7864, n_7865, n_7866, n_7867, n_7868, n_7869, n_7870;
  wire n_7871, n_7872, n_7873, n_7874, n_7875, n_7876, n_7877, n_7878;
  wire n_7879, n_7880, n_7881, n_7882, n_7883, n_7884, n_7885, n_7886;
  wire n_7887, n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894;
  wire n_7895, n_7896, n_7897, n_7898, n_7899, n_7900, n_7901, n_7902;
  wire n_7903, n_7904, n_7905, n_7906, n_7907, n_7908, n_7909, n_7910;
  wire n_7911, n_7912, n_7913, n_7914, n_7915, n_7916, n_7917, n_7918;
  wire n_7919, n_7920, n_7921, n_7922, n_7923, n_7924, n_7925, n_7926;
  wire n_7927, n_7928, n_7929, n_7930, n_7931, n_7932, n_7933, n_7934;
  wire n_7935, n_7936, n_7937, n_7938, n_7939, n_7940, n_7941, n_7942;
  wire n_7943, n_7944, n_7945, n_7946, n_7947, n_7948, n_7949, n_7950;
  wire n_7951, n_7952, n_7953, n_7954, n_7955, n_7956, n_7957, n_7958;
  wire n_7959, n_7960, n_7961, n_7962, n_7963, n_7964, n_7966, n_7967;
  wire n_7968, n_7969, n_7970, n_7971, n_7972, n_7973, n_7974, n_7975;
  wire n_7976, n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983;
  wire n_7984, n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991;
  wire n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999;
  wire n_8000, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007;
  wire n_8008, n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015;
  wire n_8016, n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023;
  wire n_8024, n_8025, n_8026, n_8027, n_8028, n_8029, n_8030, n_8031;
  wire n_8032, n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, n_8039;
  wire n_8040, n_8041, n_8042, n_8043, n_8044, n_8045, n_8046, n_8047;
  wire n_8048, n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055;
  wire n_8056, n_8057, n_8058, n_8059, n_8060, n_8061, n_8062, n_8063;
  wire n_8064, n_8065, n_8066, n_8067, n_8068, n_8069, n_8070, n_8071;
  wire n_8072, n_8073, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079;
  wire n_8080, n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087;
  wire n_8088, n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095;
  wire n_8096, n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103;
  wire n_8104, n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111;
  wire n_8112, n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8120;
  wire n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128;
  wire n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136;
  wire n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144;
  wire n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152;
  wire n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160;
  wire n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168;
  wire n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176;
  wire n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184;
  wire n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192;
  wire n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200;
  wire n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208;
  wire n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216;
  wire n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224;
  wire n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232;
  wire n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240;
  wire n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248;
  wire n_8249, n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256;
  wire n_8257, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264;
  wire n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272;
  wire n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280;
  wire n_8281, n_8282, n_8283, n_8284, n_8285, n_8286, n_8287, n_8288;
  wire n_8289, n_8290, n_8291, n_8292, n_8293, n_8294, n_8295, n_8296;
  wire n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304;
  wire n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312;
  wire n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320;
  wire n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328;
  wire n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336;
  wire n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344;
  wire n_8345, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351, n_8352;
  wire n_8353, n_8354, n_8355, n_8356, n_8357, n_8358, n_8359, n_8360;
  wire n_8361, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367, n_8368;
  wire n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376;
  wire n_8378, n_8379, n_8380, n_8381, n_8382, n_8383, n_8384, n_8385;
  wire n_8386, n_8387, n_8388, n_8389, n_8390, n_8391, n_8392, n_8393;
  wire n_8394, n_8395, n_8396, n_8397, n_8398, n_8399, n_8400, n_8401;
  wire n_8402, n_8403, n_8404, n_8405, n_8406, n_8407, n_8408, n_8409;
  wire n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416, n_8417;
  wire n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424, n_8425;
  wire n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432, n_8433;
  wire n_8434, n_8435, n_8436, n_8437, n_8438, n_8439, n_8440, n_8441;
  wire n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448, n_8449;
  wire n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456, n_8457;
  wire n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464, n_8465;
  wire n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472, n_8473;
  wire n_8474, n_8475, n_8476, n_8477, n_8478, n_8479, n_8480, n_8481;
  wire n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488, n_8489;
  wire n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496, n_8497;
  wire n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, n_8504, n_8505;
  wire n_8506, n_8507, n_8508, n_8509, n_8510, n_8511, n_8512, n_8513;
  wire n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520, n_8521;
  wire n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528, n_8529;
  wire n_8530, n_8531, n_8532, n_8533, n_8534, n_8535, n_8536, n_8537;
  wire n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544, n_8545;
  wire n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552, n_8553;
  wire n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560, n_8561;
  wire n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568, n_8569;
  wire n_8570, n_8571, n_8572, n_8573, n_8574, n_8575, n_8576, n_8577;
  wire n_8578, n_8579, n_8580, n_8581, n_8582, n_8583, n_8584, n_8585;
  wire n_8586, n_8587, n_8588, n_8589, n_8590, n_8591, n_8592, n_8593;
  wire n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600, n_8601;
  wire n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608, n_8609;
  wire n_8610, n_8611, n_8612, n_8613, n_8614, n_8615, n_8616, n_8617;
  wire n_8618, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8625;
  wire n_8626, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632, n_8633;
  wire n_8634, n_8635, n_8636, n_8637, n_8638, n_8639, n_8640, n_8641;
  wire n_8642, n_8643, n_8644, n_8645, n_8646, n_8647, n_8648, n_8649;
  wire n_8650, n_8651, n_8652, n_8653, n_8654, n_8655, n_8656, n_8657;
  wire n_8658, n_8659, n_8660, n_8661, n_8662, n_8663, n_8664, n_8665;
  wire n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, n_8672, n_8673;
  wire n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681;
  wire n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689;
  wire n_8690, n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697;
  wire n_8698, n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705;
  wire n_8706, n_8707, n_8708, n_8709, n_8710, n_8711, n_8712, n_8713;
  wire n_8714, n_8715, n_8716, n_8717, n_8718, n_8719, n_8720, n_8721;
  wire n_8722, n_8723, n_8724, n_8725, n_8726, n_8727, n_8728, n_8729;
  wire n_8730, n_8731, n_8732, n_8733, n_8734, n_8735, n_8736, n_8737;
  wire n_8738, n_8739, n_8740, n_8741, n_8742, n_8743, n_8744, n_8745;
  wire n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8752, n_8753;
  wire n_8754, n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761;
  wire n_8762, n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769;
  wire n_8770, n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777;
  wire n_8778, n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785;
  wire n_8786, n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793;
  wire n_8794, n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801;
  wire n_8802, n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8809;
  wire n_8810, n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817;
  wire n_8818, n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, n_8825;
  wire n_8826, n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833;
  wire n_8834, n_8835, n_8836, n_8837, n_8838, n_8839, n_8840, n_8841;
  wire n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8848, n_8849;
  wire n_8850, n_8851, n_8852, n_8853, n_8854, n_8855, n_8856, n_8857;
  wire n_8858, n_8859, n_8860, n_8861, n_8862, n_8863, n_8864, n_8865;
  wire n_8866, n_8867, n_8868, n_8869, n_8870, n_8871, n_8872, n_8873;
  wire n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881;
  wire n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889;
  wire n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897;
  wire n_8898, n_8899, n_8900, n_8901, n_8902, n_8903, n_8904, n_8905;
  wire n_8906, n_8907, n_8908, n_8909, n_8910, n_8911, n_8912, n_8913;
  wire n_8914, n_8915, n_8916, n_8917, n_8918, n_8919, n_8920, n_8921;
  wire n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928, n_8929;
  wire n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936, n_8937;
  wire n_8938, n_8939, n_8940, n_8941, n_8942, n_8943, n_8944, n_8945;
  wire n_8946, n_8947, n_8948, n_8949, n_8950, n_8951, n_8952, n_8953;
  wire n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960, n_8961;
  wire n_8962, n_8963, n_8964, n_8965, n_8966, n_8967, n_8968, n_8969;
  wire n_8970, n_8971, n_8972, n_8973, n_8974, n_8975, n_8976, n_8977;
  wire n_8978, n_8979, n_8980, n_8981, n_8982, n_8983, n_8984, n_8985;
  wire n_8986, n_8987, n_8988, n_8989, n_8990, n_8991, n_8992, n_8993;
  wire n_8994, n_8995, n_8996, n_8997, n_8998, n_8999, n_9000, n_9001;
  wire n_9002, n_9003, n_9004, n_9005, n_9006, n_9007, n_9008, n_9009;
  wire n_9010, n_9011, n_9012, n_9013, n_9014, n_9015, n_9016, n_9017;
  wire n_9018, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024, n_9025;
  wire n_9026, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032, n_9033;
  wire n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040, n_9041;
  wire n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048, n_9049;
  wire n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056, n_9057;
  wire n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9064, n_9065;
  wire n_9066, n_9067, n_9068, n_9069, n_9070, n_9071, n_9072, n_9073;
  wire n_9074, n_9075, n_9076, n_9077, n_9078, n_9079, n_9080, n_9081;
  wire n_9082, n_9083, n_9084, n_9085, n_9086, n_9087, n_9088, n_9089;
  wire n_9090, n_9091, n_9092, n_9093, n_9094, n_9095, n_9096, n_9097;
  wire n_9098, n_9099, n_9100, n_9101, n_9102, n_9103, n_9104, n_9105;
  wire n_9106, n_9107, n_9108, n_9109, n_9110, n_9111, n_9112, n_9113;
  wire n_9114, n_9115, n_9116, n_9117, n_9118, n_9119, n_9120, n_9121;
  wire n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128, n_9129;
  wire n_9130, n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137;
  wire n_9138, n_9139, n_9140, n_9141, n_9142, n_9143, n_9144, n_9145;
  wire n_9146, n_9147, n_9148, n_9149, n_9150, n_9151, n_9152, n_9153;
  wire n_9154, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160, n_9161;
  wire n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9168, n_9169;
  wire n_9170, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176, n_9177;
  wire n_9178, n_9179, n_9180, n_9181, n_9182, n_9183, n_9184, n_9185;
  wire n_9186, n_9187, n_9188, n_9189, n_9190, n_9191, n_9192, n_9193;
  wire n_9194, n_9195, n_9196, n_9197, n_9198, n_9199, n_9200, n_9201;
  wire n_9202, n_9203, n_9204, n_9205, n_9206, n_9207, n_9208, n_9209;
  wire n_9210, n_9211, n_9212, n_9213, n_9214, n_9215, n_9216, n_9217;
  wire n_9218, n_9219, n_9220, n_9221, n_9222, n_9223, n_9224, n_9225;
  wire n_9226, n_9227, n_9228, n_9229, n_9230, n_9231, n_9232, n_9233;
  wire n_9234, n_9235, n_9236, n_9237, n_9238, n_9239, n_9240, n_9241;
  wire n_9242, n_9243, n_9244, n_9245, n_9246, n_9247, n_9248, n_9249;
  wire n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256, n_9257;
  wire n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265;
  wire n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, n_9273;
  wire n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281;
  wire n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288, n_9289;
  wire n_9290, n_9291, n_9292, n_9293, n_9294, n_9295, n_9296, n_9297;
  wire n_9298, n_9299, n_9300, n_9301, n_9302, n_9303, n_9304, n_9305;
  wire n_9306, n_9307, n_9308, n_9309, n_9310, n_9311, n_9312, n_9313;
  wire n_9314, n_9315, n_9316, n_9317, n_9318, n_9319, n_9320, n_9321;
  wire n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9328, n_9329;
  wire n_9330, n_9331, n_9332, n_9333, n_9334, n_9335, n_9336, n_9337;
  wire n_9338, n_9339, n_9340, n_9341, n_9342, n_9343, n_9344, n_9345;
  wire n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353;
  wire n_9354, n_9355, n_9356, n_9357, n_9358, n_9359, n_9360, n_9361;
  wire n_9362, n_9363, n_9364, n_9365, n_9366, n_9367, n_9368, n_9369;
  wire n_9370, n_9371, n_9372, n_9373, n_9374, n_9375, n_9376, n_9377;
  wire n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9384, n_9385;
  wire n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, n_9392, n_9393;
  wire n_9394, n_9395, n_9396, n_9397, n_9398, n_9399, n_9400, n_9401;
  wire n_9402, n_9403, n_9404, n_9405, n_9406, n_9407, n_9408, n_9409;
  wire n_9410, n_9411, n_9412, n_9413, n_9414, n_9415, n_9416, n_9417;
  wire n_9418, n_9419, n_9420, n_9421, n_9422, n_9423, n_9424, n_9425;
  wire n_9426, n_9427, n_9428, n_9429, n_9430, n_9431, n_9432, n_9433;
  wire n_9434, n_9435, n_9436, n_9437, n_9438, n_9439, n_9440, n_9441;
  wire n_9442, n_9443, n_9444, n_9445, n_9446, n_9447, n_9448, n_9449;
  wire n_9450, n_9451, n_9452, n_9453, n_9454, n_9455, n_9456, n_9457;
  wire n_9458, n_9459, n_9460, n_9461, n_9462, n_9463, n_9464, n_9465;
  wire n_9466, n_9467, n_9468, n_9469, n_9470, n_9471, n_9472, n_9473;
  wire n_9474, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480, n_9481;
  wire n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489;
  wire n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496, n_9497;
  wire n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504, n_9505;
  wire n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512, n_9513;
  wire n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520, n_9521;
  wire n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, n_9528, n_9529;
  wire n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536, n_9537;
  wire n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545;
  wire n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552, n_9553;
  wire n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561;
  wire n_9562, n_9563, n_9564, n_9565, n_9566, n_9567, n_9568, n_9569;
  wire n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576, n_9577;
  wire n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584, n_9585;
  wire n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592, n_9593;
  wire n_9594, n_9595, n_9596, n_9597, n_9598, n_9599, n_9600, n_9601;
  wire n_9602, n_9603, n_9604, n_9605, n_9606, n_9607, n_9608, n_9609;
  wire n_9610, n_9611, n_9612, n_9613, n_9614, n_9615, n_9616, n_9617;
  wire n_9618, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624, n_9625;
  wire n_9626, n_9627, n_9628, n_9629, n_9630, n_9631, n_9632, n_9633;
  wire n_9634, n_9635, n_9636, n_9637, n_9638, n_9639, n_9640, n_9641;
  wire n_9642, n_9643, n_9644, n_9645, n_9646, n_9647, n_9648, n_9649;
  wire n_9650, n_9651, n_9652, n_9653, n_9654, n_9655, n_9656, n_9657;
  wire n_9658, n_9659, n_9660, n_9661, n_9662, n_9663, n_9664, n_9665;
  wire n_9666, n_9667, n_9668, n_9669, n_9670, n_9671, n_9672, n_9673;
  wire n_9674, n_9675, n_9676, n_9677, n_9678, n_9679, n_9680, n_9681;
  wire n_9682, n_9683, n_9684, n_9685, n_9686, n_9687, n_9688, n_9689;
  wire n_9690, n_9691, n_9692, n_9693, n_9694, n_9695, n_9696, n_9697;
  wire n_9698, n_9699, n_9700, n_9701, n_9702, n_9703, n_9704, n_9705;
  wire n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712, n_9713;
  wire n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720, n_9721;
  wire n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728, n_9729;
  wire n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736, n_9737;
  wire n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744, n_9745;
  wire n_9746, n_9747, n_9748, n_9749, n_9750, n_9751, n_9752, n_9753;
  wire n_9754, n_9755, n_9756, n_9757, n_9758, n_9759, n_9760, n_9761;
  wire n_9762, n_9763, n_9764, n_9765, n_9766, n_9767, n_9768, n_9769;
  wire n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776, n_9777;
  wire n_9778, n_9779, n_9780, n_9781, n_9782, n_9783, n_9784, n_9785;
  wire n_9786, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792, n_9793;
  wire n_9794, n_9795, n_9796, n_9797, n_9798, n_9799, n_9800, n_9801;
  wire n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808, n_9809;
  wire n_9810, n_9811, n_9812, n_9813, n_9814, n_9815, n_9816, n_9817;
  wire n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_9825;
  wire n_9826, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832, n_9833;
  wire n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841;
  wire n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848, n_9849;
  wire n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856, n_9857;
  wire n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864, n_9865;
  wire n_9866, n_9867, n_9868, n_9869, n_9870, n_9871, n_9872, n_9873;
  wire n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880, n_9881;
  wire n_9882, n_9883, n_9884, n_9885, n_9886, n_9887, n_9888, n_9889;
  wire n_9890, n_9891, n_9892, n_9893, n_9894, n_9895, n_9896, n_9897;
  wire n_9898, n_9899, n_9900, n_9901, n_9902, n_9903, n_9904, n_9905;
  wire n_9906, n_9907, n_9908, n_9909, n_9910, n_9911, n_9912, n_9913;
  wire n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920, n_9921;
  wire n_9922, n_9923, n_9924, n_9925, n_9926, n_9927, n_9928, n_9929;
  wire n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937;
  wire n_9938, n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945;
  wire n_9946, n_9947, n_9948, n_9949, n_9950, n_9951, n_9952, n_9953;
  wire n_9954, n_9955, n_9956, n_9957, n_9958, n_9959, n_9960, n_9961;
  wire n_9962, n_9963, n_9964, n_9965, n_9966, n_9967, n_9968, n_9969;
  wire n_9970, n_9971, n_9972, n_9973, n_9974, n_9975, n_9976, n_9977;
  wire n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984, n_9985;
  wire n_9986, n_9987, n_9988, n_9989, n_9990, n_9991, n_9992, n_9993;
  wire n_9994, n_9995, n_9996, n_9997, n_9998, n_9999, n_10000, n_10001;
  wire n_10002, n_10003, n_10004, n_10005, n_10006, n_10007, n_10008,
       n_10009;
  wire n_10010, n_10011, n_10012, n_10013, n_10014, n_10015, n_10016,
       n_10017;
  wire n_10018, n_10019, n_10020, n_10021, n_10022, n_10023, n_10024,
       n_10025;
  wire n_10026, n_10027, n_10028, n_10029, n_10030, n_10031, n_10032,
       n_10033;
  wire n_10034, n_10035, n_10036, n_10037, n_10038, n_10039, n_10040,
       n_10041;
  wire n_10042, n_10043, n_10044, n_10045, n_10046, n_10047, n_10048,
       n_10049;
  wire n_10050, n_10051, n_10052, n_10053, n_10054, n_10055, n_10056,
       n_10057;
  wire n_10058, n_10059, n_10060, n_10061, n_10062, n_10063, n_10064,
       n_10065;
  wire n_10066, n_10067, n_10068, n_10069, n_10070, n_10071, n_10072,
       n_10073;
  wire n_10074, n_10075, n_10076, n_10077, n_10078, n_10079, n_10080,
       n_10081;
  wire n_10082, n_10083, n_10084, n_10085, n_10086, n_10087, n_10088,
       n_10089;
  wire n_10090, n_10091, n_10092, n_10093, n_10094, n_10095, n_10096,
       n_10097;
  wire n_10098, n_10099, n_10100, n_10101, n_10102, n_10103, n_10104,
       n_10105;
  wire n_10106, n_10107, n_10108, n_10109, n_10110, n_10111, n_10112,
       n_10113;
  wire n_10114, n_10115, n_10116, n_10117, n_10118, n_10119, n_10120,
       n_10121;
  wire n_10122, n_10123, n_10124, n_10125, n_10126, n_10127, n_10128,
       n_10129;
  wire n_10130, n_10131, n_10132, n_10133, n_10134, n_10135, n_10136,
       n_10137;
  wire n_10138, n_10139, n_10140, n_10141, n_10142, n_10143, n_10144,
       n_10145;
  wire n_10146, n_10147, n_10148, n_10149, n_10150, n_10151, n_10152,
       n_10153;
  wire n_10154, n_10155, n_10156, n_10157, n_10158, n_10159, n_10160,
       n_10161;
  wire n_10162, n_10163, n_10164, n_10165, n_10166, n_10167, n_10168,
       n_10169;
  wire n_10170, n_10171, n_10172, n_10173, n_10174, n_10175, n_10176,
       n_10177;
  wire n_10178, n_10179, n_10180, n_10181, n_10182, n_10183, n_10184,
       n_10185;
  wire n_10186, n_10187, n_10188, n_10189, n_10190, n_10191, n_10192,
       n_10193;
  wire n_10194, n_10195, n_10196, n_10197, n_10198, n_10199, n_10200,
       n_10201;
  wire n_10202, n_10203, n_10204, n_10205, n_10206, n_10207, n_10208,
       n_10209;
  wire n_10210, n_10211, n_10212, n_10213, n_10214, n_10215, n_10216,
       n_10217;
  wire n_10218, n_10219, n_10220, n_10221, n_10222, n_10223, n_10224,
       n_10225;
  wire n_10226, n_10227, n_10228, n_10229, n_10230, n_10231, n_10232,
       n_10233;
  wire n_10234, n_10235, n_10236, n_10237, n_10238, n_10239, n_10240,
       n_10241;
  wire n_10242, n_10243, n_10244, n_10245, n_10246, n_10247, n_10248,
       n_10249;
  wire n_10250, n_10251, n_10252, n_10253, n_10254, n_10255, n_10256,
       n_10257;
  wire n_10258, n_10259, n_10260, n_10261, n_10262, n_10263, n_10264,
       n_10265;
  wire n_10266, n_10267, n_10268, n_10269, n_10270, n_10271, n_10272,
       n_10273;
  wire n_10274, n_10275, n_10276, n_10277, n_10278, n_10279, n_10280,
       n_10281;
  wire n_10282, n_10283, n_10284, n_10285, n_10286, n_10287, n_10288,
       n_10289;
  wire n_10290, n_10291, n_10292, n_10293, n_10294, n_10295, n_10296,
       n_10297;
  wire n_10298, n_10299, n_10300, n_10301, n_10302, n_10303, n_10304,
       n_10305;
  wire n_10306, n_10307, n_10308, n_10309, n_10310, n_10311, n_10312,
       n_10313;
  wire n_10314, n_10315, n_10316, n_10317, n_10318, n_10319, n_10320,
       n_10321;
  wire n_10322, n_10323, n_10324, n_10325, n_10326, n_10327, n_10328,
       n_10329;
  wire n_10330, n_10331, n_10332, n_10333, n_10334, n_10335, n_10336,
       n_10337;
  wire n_10338, n_10339, n_10340, n_10341, n_10342, n_10343, n_10344,
       n_10345;
  wire n_10346, n_10347, n_10348, n_10349, n_10350, n_10351, n_10352,
       n_10353;
  wire n_10354, n_10355, n_10356, n_10357, n_10358, n_10359, n_10360,
       n_10361;
  wire n_10362, n_10363, n_10364, n_10365, n_10366, n_10367, n_10368,
       n_10369;
  wire n_10370, n_10371, n_10372, n_10373, n_10374, n_10375, n_10376,
       n_10377;
  wire n_10378, n_10379, n_10380, n_10381, n_10382, n_10383, n_10384,
       n_10385;
  wire n_10386, n_10387, n_10388, n_10389, n_10390, n_10391, n_10392,
       n_10393;
  wire n_10394, n_10395, n_10396, n_10397, n_10398, n_10399, n_10400,
       n_10401;
  wire n_10402, n_10403, n_10404, n_10405, n_10406, n_10407, n_10408,
       n_10409;
  wire n_10410, n_10411, n_10412, n_10413, n_10414, n_10415, n_10416,
       n_10417;
  wire n_10418, n_10419, n_10420, n_10421, n_10422, n_10423, n_10424,
       n_10425;
  wire n_10426, n_10427, n_10428, n_10429, n_10430, n_10431, n_10432,
       n_10433;
  wire n_10434, n_10435, n_10436, n_10437, n_10438, n_10439, n_10440,
       n_10441;
  wire n_10442, n_10443, n_10444, n_10445, n_10446, n_10447, n_10448,
       n_10449;
  wire n_10450, n_10451, n_10452, n_10453, n_10454, n_10455, n_10456,
       n_10457;
  wire n_10458, n_10459, n_10460, n_10461, n_10462, n_10463, n_10464,
       n_10465;
  wire n_10466, n_10467, n_10468, n_10469, n_10470, n_10471, n_10472,
       n_10473;
  wire n_10474, n_10475, n_10476, n_10477, n_10478, n_10479, n_10480,
       n_10481;
  wire n_10482, n_10483, n_10484, n_10485, n_10486, n_10487, n_10488,
       n_10489;
  wire n_10490, n_10491, n_10492, n_10493, n_10494, n_10495, n_10496,
       n_10497;
  wire n_10498, n_10499, n_10500, n_10501, n_10502, n_10503, n_10504,
       n_10505;
  wire n_10506, n_10507, n_10508, n_10509, n_10510, n_10511, n_10512,
       n_10513;
  wire n_10514, n_10515, n_10516, n_10517, n_10518, n_10519, n_10520,
       n_10521;
  wire n_10522, n_10523, n_10524, n_10525, n_10526, n_10527, n_10528,
       n_10529;
  wire n_10530, n_10531, n_10532, n_10533, n_10534, n_10535, n_10536,
       n_10537;
  wire n_10538, n_10539, n_10540, n_10541, n_10542, n_10543, n_10544,
       n_10545;
  wire n_10546, n_10547, n_10548, n_10549, n_10550, n_10551, n_10552,
       n_10553;
  wire n_10554, n_10555, n_10556, n_10557, n_10558, n_10559, n_10560,
       n_10561;
  wire n_10562, n_10563, n_10564, n_10565, n_10566, n_10567, n_10568,
       n_10569;
  wire n_10570, n_10571, n_10572, n_10573, n_10574, n_10575, n_10576,
       n_10577;
  wire n_10578, n_10579, n_10580, n_10581, n_10582, n_10583, n_10584,
       n_10585;
  wire n_10586, n_10587, n_10588, n_10589, n_10590, n_10591, n_10592,
       n_10593;
  wire n_10594, n_10595, n_10596, n_10597, n_10598, n_10599, n_10600,
       n_10601;
  wire n_10602, n_10603, n_10604, n_10605, n_10606, n_10607, n_10608,
       n_10609;
  wire n_10610, n_10611, n_10612, n_10613, n_10614, n_10615, n_10616,
       n_10617;
  wire n_10618, n_10619, n_10620, n_10621, n_10622, n_10623, n_10624,
       n_10625;
  wire n_10626, n_10627, n_10628, n_10629, n_10630, n_10631, n_10632,
       n_10633;
  wire n_10634, n_10635, n_10636, n_10637, n_10638, n_10639, n_10640,
       n_10641;
  wire n_10642, n_10643, n_10644, n_10645, n_10646, n_10647, n_10648,
       n_10649;
  wire n_10650, n_10651, n_10652, n_10653, n_10654, n_10655, n_10656,
       n_10657;
  wire n_10658, n_10659, n_10660, n_10661, n_10662, n_10663, n_10664,
       n_10665;
  wire n_10666, n_10667, n_10668, n_10669, n_10670, n_10671, n_10672,
       n_10673;
  wire n_10674, n_10675, n_10676, n_10677, n_10678, n_10679, n_10680,
       n_10681;
  wire n_10682, n_10683, n_10684, n_10685, n_10686, n_10687, n_10688,
       n_10689;
  wire n_10690, n_10691, n_10692, n_10693, n_10694, n_10695, n_10696,
       n_10697;
  wire n_10698, n_10699, n_10700, n_10701, n_10702, n_10703, n_10704,
       n_10705;
  wire n_10706, n_10707, n_10708, n_10709, n_10710, n_10711, n_10712,
       n_10713;
  wire n_10714, n_10715, n_10716, n_10717, n_10718, n_10719, n_10720,
       n_10721;
  wire n_10722, n_10723, n_10724, n_10725, n_10726, n_10727, n_10728,
       n_10729;
  wire n_10730, n_10731, n_10732, n_10733, n_10734, n_10735, n_10736,
       n_10737;
  wire n_10738, n_10739, n_10740, n_10741, n_10742, n_10743, n_10744,
       n_10745;
  wire n_10746, n_10747, n_10748, n_10749, n_10750, n_10751, n_10752,
       n_10753;
  wire n_10754, n_10755, n_10756, n_10757, n_10758, n_10759, n_10760,
       n_10761;
  wire n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768,
       n_10769;
  wire n_10770, n_10771, n_10772, n_10773, n_10774, n_10775, n_10776,
       n_10777;
  wire n_10778, n_10779, n_10780, n_10781, n_10782, n_10783, n_10784,
       n_10785;
  wire n_10786, n_10787, n_10788, n_10789, n_10790, n_10791, n_10792,
       n_10793;
  wire n_10794, n_10795, n_10796, n_10797, n_10798, n_10799, n_10800,
       n_10801;
  wire n_10802, n_10803, n_10804, n_10805, n_10806, n_10807, n_10808,
       n_10809;
  wire n_10810, n_10811, n_10812, n_10813, n_10814, n_10815, n_10816,
       n_10817;
  wire n_10818, n_10819, n_10820, n_10821, n_10822, n_10823, n_10824,
       n_10825;
  wire n_10826, n_10827, n_10828, n_10829, n_10830, n_10831, n_10832,
       n_10833;
  wire n_10834, n_10835, n_10836, n_10837, n_10838, n_10839, n_10840,
       n_10841;
  wire n_10842, n_10843, n_10844, n_10845, n_10846, n_10847, n_10848,
       n_10849;
  wire n_10850, n_10851, n_10852, n_10853, n_10854, n_10855, n_10856,
       n_10857;
  wire n_10858, n_10859, n_10860, n_10861, n_10862, n_10863, n_10864,
       n_10865;
  wire n_10866, n_10867, n_10868, n_10869, n_10870, n_10871, n_10872,
       n_10873;
  wire n_10874, n_10875, n_10876, n_10877, n_10878, n_10879, n_10880,
       n_10881;
  wire n_10882, n_10883, n_10884, n_10885, n_10886, n_10887, n_10888,
       n_10889;
  wire n_10890, n_10891, n_10892, n_10893, n_10894, n_10895, n_10896,
       n_10897;
  wire n_10898, n_10899, n_10900, n_10901, n_10902, n_10903, n_10904,
       n_10905;
  wire n_10906, n_10907, n_10908, n_10909, n_10910, n_10911, n_10912,
       n_10913;
  wire n_10914, n_10915, n_10916, n_10917, n_10918, n_10919, n_10920,
       n_10921;
  wire n_10922, n_10923, n_10924, n_10925, n_10926, n_10927, n_10928,
       n_10929;
  wire n_10930, n_10931, n_10932, n_10933, n_10934, n_10935, n_10936,
       n_10937;
  wire n_10938, n_10939, n_10940, n_10941, n_10942, n_10943, n_10944,
       n_10945;
  wire n_10946, n_10947, n_10948, n_10949, n_10950, n_10951, n_10952,
       n_10953;
  wire n_10954, n_10955, n_10956, n_10957, n_10958, n_10959, n_10960,
       n_10961;
  wire n_10962, n_10963, n_10964, n_10965, n_10966, n_10967, n_10968,
       n_10969;
  wire n_10970, n_10971, n_10972, n_10973, n_10974, n_10975, n_10976,
       n_10977;
  wire n_10978, n_10979, n_10980, n_10981, n_10982, n_10983, n_10984,
       n_10985;
  wire n_10986, n_10987, n_10988, n_10989, n_10990, n_10991, n_10992,
       n_10993;
  wire n_10994, n_10995, n_10996, n_10997, n_10998, n_10999, n_11000,
       n_11001;
  wire n_11002, n_11003, n_11004, n_11005, n_11006, n_11007, n_11008,
       n_11009;
  wire n_11010, n_11011, n_11012, n_11013, n_11014, n_11015, n_11016,
       n_11017;
  wire n_11018, n_11019, n_11020, n_11021, n_11022, n_11023, n_11024,
       n_11025;
  wire n_11026, n_11027, n_11028, n_11029, n_11030, n_11031, n_11032,
       n_11033;
  wire n_11034, n_11035, n_11036, n_11037, n_11038, n_11039, n_11040,
       n_11041;
  wire n_11042, n_11043, n_11044, n_11045, n_11046, n_11047, n_11048,
       n_11049;
  wire n_11050, n_11051, n_11052, n_11053, n_11054, n_11055, n_11056,
       n_11057;
  wire n_11058, n_11059, n_11060, n_11061, n_11062, n_11063, n_11064,
       n_11065;
  wire n_11066, n_11067, n_11068, n_11069, n_11070, n_11071, n_11072,
       n_11073;
  wire n_11074, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080,
       n_11081;
  wire n_11082, n_11083, n_11084, n_11085, n_11086, n_11087, n_11088,
       n_11089;
  wire n_11090, n_11091, n_11092, n_11093, n_11094, n_11095, n_11096,
       n_11097;
  wire n_11098, n_11099, n_11100, n_11101, n_11102, n_11103, n_11104,
       n_11105;
  wire n_11106, n_11107, n_11108, n_11109, n_11110, n_11111, n_11112,
       n_11113;
  wire n_11114, n_11115, n_11116, n_11117, n_11118, n_11119, n_11120,
       n_11121;
  wire n_11122, n_11123, n_11124, n_11125, n_11126, n_11127, n_11128,
       n_11129;
  wire n_11130, n_11131, n_11132, n_11133, n_11134, n_11135, n_11136,
       n_11137;
  wire n_11138, n_11139, n_11140, n_11141, n_11142, n_11143, n_11144,
       n_11145;
  wire n_11146, n_11147, n_11148, n_11149, n_11150, n_11151, n_11152,
       n_11153;
  wire n_11154, n_11155, n_11156, n_11157, n_11158, n_11159, n_11160,
       n_11161;
  wire n_11162, n_11163, n_11164, n_11165, n_11166, n_11167, n_11168,
       n_11169;
  wire n_11170, n_11171, n_11172, n_11173, n_11174, n_11175, n_11176,
       n_11177;
  wire n_11178, n_11179, n_11180, n_11181, n_11182, n_11183, n_11184,
       n_11185;
  wire n_11186, n_11187, n_11188, n_11189, n_11190, n_11191, n_11192,
       n_11193;
  wire n_11194, n_11195, n_11196, n_11197, n_11198, n_11199, n_11200,
       n_11201;
  wire n_11202, n_11203, n_11204, n_11205, n_11206, n_11207, n_11208,
       n_11209;
  wire n_11210, n_11211, n_11212, n_11213, n_11214, n_11215, n_11216,
       n_11217;
  wire n_11218, n_11219, n_11220, n_11221, n_11222, n_11223, n_11224,
       n_11225;
  wire n_11226, n_11227, n_11228, n_11229, n_11230, n_11231, n_11232,
       n_11233;
  wire n_11234, n_11235, n_11236, n_11237, n_11238, n_11239, n_11240,
       n_11241;
  wire n_11242, n_11243, n_11244, n_11245, n_11246, n_11247, n_11248,
       n_11249;
  wire n_11250, n_11251, n_11252, n_11253, n_11254, n_11255, n_11256,
       n_11257;
  wire n_11258, n_11259, n_11260, n_11261, n_11262, n_11263, n_11264,
       n_11265;
  wire n_11266, n_11267, n_11268, n_11269, n_11270, n_11271, n_11272,
       n_11273;
  wire n_11274, n_11275, n_11276, n_11277, n_11278, n_11279, n_11280,
       n_11281;
  wire n_11282, n_11283, n_11284, n_11285, n_11286, n_11287, n_11288,
       n_11289;
  wire n_11290, n_11291, n_11292, n_11293, n_11294, n_11295, n_11296,
       n_11297;
  wire n_11298, n_11299, n_11300, n_11301, n_11302, n_11303, n_11304,
       n_11305;
  wire n_11306, n_11307, n_11308, n_11309, n_11310, n_11311, n_11312,
       n_11313;
  wire n_11314, n_11315, n_11316, n_11317, n_11318, n_11319, n_11320,
       n_11321;
  wire n_11322, n_11323, n_11324, n_11325, n_11326, n_11327, n_11328,
       n_11329;
  wire n_11330, n_11331, n_11332, n_11333, n_11334, n_11335, n_11336,
       n_11337;
  wire n_11338, n_11339, n_11340, n_11341, n_11342, n_11343, n_11344,
       n_11345;
  wire n_11346, n_11347, n_11348, n_11349, n_11350, n_11351, n_11352,
       n_11353;
  wire n_11354, n_11355, n_11356, n_11357, n_11358, n_11359, n_11360,
       n_11361;
  wire n_11362, n_11363, n_11364, n_11365, n_11366, n_11367, n_11368,
       n_11369;
  wire n_11370, n_11371, n_11372, n_11373, n_11374, n_11375, n_11376,
       n_11377;
  wire n_11378, n_11379, n_11380, n_11381, n_11382, n_11383, n_11384,
       n_11385;
  wire n_11386, n_11387, n_11388, n_11389, n_11390, n_11391, n_11392,
       n_11393;
  wire n_11394, n_11395, n_11396, n_11397, n_11398, n_11399, n_11400,
       n_11401;
  wire n_11402, n_11403, n_11404, n_11405, n_11406, n_11407, n_11408,
       n_11409;
  wire n_11410, n_11411, n_11412, n_11413, n_11414, n_11415, n_11416,
       n_11417;
  wire n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424,
       n_11425;
  wire n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432,
       n_11433;
  wire n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440,
       n_11441;
  wire n_11442, n_11443, n_11444, n_11445, n_11446, n_11447, n_11448,
       n_11449;
  wire n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11456,
       n_11457;
  wire n_11458, n_11459, n_11460, n_11461, n_11462, n_11463, n_11464,
       n_11465;
  wire n_11466, n_11467, n_11468, n_11469, n_11470, n_11471, n_11472,
       n_11473;
  wire n_11474, n_11475, n_11476, n_11477, n_11478, n_11479, n_11480,
       n_11481;
  wire n_11482, n_11483, n_11484, n_11485, n_11486, n_11487, n_11488,
       n_11489;
  wire n_11490, n_11491, n_11492, n_11493, n_11494, n_11495, n_11496,
       n_11497;
  wire n_11498, n_11499, n_11500, n_11501, n_11502, n_11503, n_11504,
       n_11505;
  wire n_11506, n_11507, n_11508, n_11509, n_11510, n_11511, n_11512,
       n_11513;
  wire n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520,
       n_11521;
  wire n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528,
       n_11529;
  wire n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536,
       n_11537;
  wire n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544,
       n_11545;
  wire n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552,
       n_11553;
  wire n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560,
       n_11561;
  wire n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568,
       n_11569;
  wire n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576,
       n_11577;
  wire n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584,
       n_11585;
  wire n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592,
       n_11593;
  wire n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600,
       n_11601;
  wire n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11608,
       n_11609;
  wire n_11610, n_11611, n_11612, n_11613, n_11614, n_11615, n_11616,
       n_11617;
  wire n_11618, n_11619, n_11620, n_11621, n_11622, n_11623, n_11624,
       n_11625;
  wire n_11626, n_11627, n_11628, n_11629, n_11630, n_11631, n_11632,
       n_11633;
  wire n_11634, n_11635, n_11636, n_11637, n_11638, n_11639, n_11640,
       n_11641;
  wire n_11642, n_11643, n_11644, n_11645, n_11646, n_11647, n_11648,
       n_11649;
  wire n_11650, n_11651, n_11652, n_11653, n_11654, n_11655, n_11656,
       n_11657;
  wire n_11658, n_11659, n_11660, n_11661, n_11662, n_11663, n_11664,
       n_11665;
  wire n_11666, n_11667, n_11668, n_11669, n_11670, n_11671, n_11672,
       n_11673;
  wire n_11674, n_11675, n_11676, n_11677, n_11678, n_11679, n_11680,
       n_11681;
  wire n_11682, n_11683, n_11684, n_11685, n_11686, n_11687, n_11688,
       n_11689;
  wire n_11690, n_11691, n_11692, n_11693, n_11694, n_11695, n_11696,
       n_11697;
  wire n_11698, n_11699, n_11700, n_11701, n_11702, n_11703, n_11704,
       n_11705;
  wire n_11706, n_11707, n_11708, n_11709, n_11710, n_11711, n_11712,
       n_11713;
  wire n_11714, n_11715, n_11716, n_11717, n_11718, n_11719, n_11720,
       n_11721;
  wire n_11722, n_11723, n_11724, n_11725, n_11726, n_11727, n_11728,
       n_11729;
  wire n_11730, n_11731, n_11732, n_11733, n_11734, n_11735, n_11736,
       n_11737;
  wire n_11738, n_11739, n_11740, n_11741, n_11742, n_11743, n_11744,
       n_11745;
  wire n_11746, n_11747, n_11748, n_11749, n_11750, n_11751, n_11752,
       n_11753;
  wire n_11754, n_11755, n_11756, n_11757, n_11758, n_11759, n_11760,
       n_11761;
  wire n_11762, n_11763, n_11764, n_11765, n_11766, n_11767, n_11768,
       n_11769;
  wire n_11770, n_11771, n_11772, n_11773, n_11774, n_11775, n_11776,
       n_11777;
  wire n_11778, n_11779, n_11780, n_11781, n_11782, n_11783, n_11784,
       n_11785;
  wire n_11786, n_11787, n_11788, n_11789, n_11790, n_11791, n_11792,
       n_11793;
  wire n_11794, n_11795, n_11796, n_11797, n_11798, n_11799, n_11800,
       n_11801;
  wire n_11802, n_11803, n_11804, n_11805, n_11806, n_11807, n_11808,
       n_11809;
  wire n_11810, n_11811, n_11812, n_11813, n_11814, n_11815, n_11816,
       n_11817;
  wire n_11818, n_11819, n_11820, n_11821, n_11822, n_11823, n_11824,
       n_11825;
  wire n_11826, n_11827, n_11828, n_11829, n_11830, n_11831, n_11832,
       n_11833;
  wire n_11834, n_11835, n_11836, n_11837, n_11838, n_11839, n_11840,
       n_11841;
  wire n_11842, n_11843, n_11844, n_11845, n_11846, n_11847, n_11848,
       n_11849;
  wire n_11850, n_11851, n_11852, n_11853, n_11854, n_11855, n_11856,
       n_11857;
  wire n_11858, n_11859, n_11860, n_11861, n_11862, n_11863, n_11864,
       n_11865;
  wire n_11866, n_11867, n_11868, n_11869, n_11870, n_11871, n_11872,
       n_11873;
  wire n_11874, n_11875, n_11876, n_11877, n_11878, n_11879, n_11880,
       n_11881;
  wire n_11882, n_11883, n_11884, n_11885, n_11886, n_11887, n_11888,
       n_11889;
  wire n_11890, n_11891, n_11892, n_11893, n_11894, n_11895, n_11896,
       n_11897;
  wire n_11898, n_11899, n_11900, n_11901, n_11902, n_11903, n_11904,
       n_11905;
  wire n_11906, n_11907, n_11908, n_11909, n_11910, n_11911, n_11912,
       n_11913;
  wire n_11914, n_11915, n_11916, n_11917, n_11918, n_11919, n_11920,
       n_11921;
  wire n_11922, n_11923, n_11924, n_11925, n_11926, n_11927, n_11928,
       n_11929;
  wire n_11930, n_11931, n_11932, n_11933, n_11934, n_11935, n_11936,
       n_11937;
  wire n_11938, n_11939, n_11940, n_11941, n_11942, n_11943, n_11944,
       n_11945;
  wire n_11946, n_11947, n_11948, n_11949, n_11950, n_11951, n_11952,
       n_11953;
  wire n_11954, n_11955, n_11956, n_11957, n_11958, n_11959, n_11960,
       n_11961;
  wire n_11962, n_11963, n_11964, n_11965, n_11966, n_11967, n_11968,
       n_11969;
  wire n_11970, n_11971, n_11972, n_11973, n_11974, n_11975, n_11976,
       n_11977;
  wire n_11978, n_11979, n_11980, n_11981, n_11982, n_11983, n_11984,
       n_11985;
  wire n_11986, n_11987, n_11988, n_11989, n_11990, n_11991, n_11992,
       n_11993;
  wire n_11994, n_11995, n_11996, n_11997, n_11998, n_11999, n_12000,
       n_12001;
  wire n_12002, n_12003, n_12004, n_12005, n_12006, n_12007, n_12008,
       n_12009;
  wire n_12010, n_12011, n_12012, n_12013, n_12014, n_12015, n_12016,
       n_12017;
  wire n_12018, n_12019, n_12020, n_12021, n_12022, n_12023, n_12024,
       n_12025;
  wire n_12026, n_12027, n_12028, n_12029, n_12030, n_12031, n_12032,
       n_12033;
  wire n_12034, n_12035, n_12036, n_12037, n_12038, n_12039, n_12040,
       n_12041;
  wire n_12042, n_12043, n_12044, n_12045, n_12046, n_12047, n_12048,
       n_12049;
  wire n_12050, n_12051, n_12052, n_12053, n_12054, n_12055, n_12056,
       n_12057;
  wire n_12058, n_12059, n_12060, n_12061, n_12062, n_12063, n_12064,
       n_12065;
  wire n_12066, n_12067, n_12068, n_12069, n_12070, n_12071, n_12072,
       n_12073;
  wire n_12074, n_12075, n_12076, n_12077, n_12078, n_12079, n_12080,
       n_12081;
  wire n_12082, n_12083, n_12084, n_12085, n_12086, n_12087, n_12088,
       n_12089;
  wire n_12090, n_12091, n_12092, n_12093, n_12094, n_12095, n_12096,
       n_12097;
  wire n_12098, n_12099, n_12100, n_12101, n_12102, n_12103, n_12104,
       n_12105;
  wire n_12106, n_12107, n_12108, n_12109, n_12110, n_12111, n_12112,
       n_12113;
  wire n_12114, n_12115, n_12116, n_12117, n_12118, n_12119, n_12120,
       n_12121;
  wire n_12122, n_12123, n_12124, n_12125, n_12126, n_12127, n_12128,
       n_12129;
  wire n_12130, n_12131, n_12132, n_12133, n_12134, n_12135, n_12136,
       n_12137;
  wire n_12138, n_12139, n_12140, n_12141, n_12142, n_12143, n_12144,
       n_12145;
  wire n_12146, n_12147, n_12148, n_12149, n_12150, n_12151, n_12152,
       n_12153;
  wire n_12154, n_12155, n_12156, n_12157, n_12158, n_12159, n_12160,
       n_12161;
  wire n_12162, n_12163, n_12164, n_12165, n_12166, n_12167, n_12168,
       n_12169;
  wire n_12170, n_12171, n_12172, n_12173, n_12174, n_12175, n_12176,
       n_12177;
  wire n_12178, n_12179, n_12180, n_12181, n_12182, n_12183, n_12184,
       n_12185;
  wire n_12186, n_12187, n_12188, n_12189, n_12190, n_12191, n_12192,
       n_12193;
  wire n_12194, n_12195, n_12196, n_12197, n_12198, n_12199, n_12200,
       n_12201;
  wire n_12202, n_12203, n_12204, n_12205, n_12206, n_12207, n_12208,
       n_12209;
  wire n_12210, n_12211, n_12212, n_12213, n_12214, n_12215, n_12216,
       n_12217;
  wire n_12218, n_12219, n_12220, n_12221, n_12222, n_12223, n_12224,
       n_12225;
  wire n_12226, n_12227, n_12228, n_12229, n_12230, n_12231, n_12232,
       n_12233;
  wire n_12234, n_12235, n_12236, n_12237, n_12238, n_12239, n_12240,
       n_12241;
  wire n_12242, n_12243, n_12244, n_12245, n_12246, n_12247, n_12248,
       n_12249;
  wire n_12250, n_12251, n_12252, n_12253, n_12254, n_12255, n_12256,
       n_12257;
  wire n_12258, n_12259, n_12260, n_12261, n_12262, n_12263, n_12264,
       n_12265;
  wire n_12266, n_12267, n_12268, n_12269, n_12270, n_12271, n_12272,
       n_12273;
  wire n_12274, n_12275, n_12276, n_12277, n_12278, n_12279, n_12280,
       n_12281;
  wire n_12282, n_12283, n_12284, n_12285, n_12286, n_12287, n_12288,
       n_12289;
  wire n_12290, n_12291, n_12292, n_12293, n_12294, n_12295, n_12296,
       n_12297;
  wire n_12298, n_12299, n_12300, n_12301, n_12302, n_12303, n_12304,
       n_12305;
  wire n_12306, n_12307, n_12308, n_12309, n_12310, n_12311, n_12312,
       n_12313;
  wire n_12314, n_12315, n_12316, n_12317, n_12318, n_12319, n_12320,
       n_12321;
  wire n_12322, n_12323, n_12324, n_12325, n_12326, n_12327, n_12328,
       n_12329;
  wire n_12330, n_12331, n_12332, n_12333, n_12334, n_12335, n_12336,
       n_12337;
  wire n_12338, n_12339, n_12340, n_12341, n_12342, n_12343, n_12344,
       n_12345;
  wire n_12346, n_12347, n_12348, n_12349, n_12350, n_12351, n_12352,
       n_12353;
  wire n_12354, n_12355, n_12356, n_12357, n_12358, n_12359, n_12360,
       n_12361;
  wire n_12362, n_12363, n_12364, n_12365, n_12366, n_12367, n_12368,
       n_12369;
  wire n_12370, n_12371, n_12372, n_12373, n_12374, n_12375, n_12376,
       n_12377;
  wire n_12378, n_12379, n_12380, n_12381, n_12382, n_12383, n_12384,
       n_12385;
  wire n_12386, n_12387, n_12388, n_12389, n_12390, n_12391, n_12392,
       n_12393;
  wire n_12394, n_12395, n_12396, n_12397, n_12398, n_12399, n_12400,
       n_12401;
  wire n_12402, n_12403, n_12404, n_12405, n_12406, n_12407, n_12408,
       n_12409;
  wire n_12410, n_12411, n_12412, n_12413, n_12414, n_12415, n_12416,
       n_12417;
  wire n_12418, n_12419, n_12420, n_12421, n_12422, n_12423, n_12424,
       n_12425;
  wire n_12426, n_12427, n_12428, n_12429, n_12430, n_12431, n_12432,
       n_12433;
  wire n_12434, n_12435, n_12436, n_12437, n_12438, n_12439, n_12440,
       n_12441;
  wire n_12442, n_12443, n_12444, n_12445, n_12446, n_12447, n_12448,
       n_12449;
  wire n_12450, n_12451, n_12452, n_12453, n_12454, n_12455, n_12456,
       n_12457;
  wire n_12458, n_12459, n_12460, n_12461, n_12462, n_12463, n_12464,
       n_12465;
  wire n_12466, n_12467, n_12468, n_12469, n_12470, n_12471, n_12472,
       n_12473;
  wire n_12474, n_12475, n_12476, n_12477, n_12478, n_12479, n_12480,
       n_12481;
  wire n_12482, n_12483, n_12484, n_12485, n_12486, n_12487, n_12488,
       n_12489;
  wire n_12490, n_12491, n_12492, n_12493, n_12494, n_12495, n_12496,
       n_12497;
  wire n_12498, n_12499, n_12500, n_12501, n_12502, n_12503, n_12504,
       n_12505;
  wire n_12506, n_12507, n_12508, n_12509, n_12510, n_12511, n_12512,
       n_12513;
  wire n_12514, n_12515, n_12516, n_12517, n_12518, n_12519, n_12520,
       n_12521;
  wire n_12522, n_12523, n_12524, n_12525, n_12526, n_12527, n_12528,
       n_12529;
  wire n_12530, n_12531, n_12532, n_12533, n_12534, n_12535, n_12536,
       n_12537;
  wire n_12538, n_12539, n_12540, n_12541, n_12542, n_12543, n_12544,
       n_12545;
  wire n_12546, n_12547, n_12548, n_12549, n_12550, n_12551, n_12552,
       n_12553;
  wire n_12554, n_12555, n_12556, n_12557, n_12558, n_12559, n_12560,
       n_12561;
  wire n_12562, n_12563, n_12564, n_12565, n_12566, n_12567, n_12568,
       n_12569;
  wire n_12570, n_12571, n_12572, n_12573, n_12574, n_12575, n_12576,
       n_12577;
  wire n_12578, n_12579, n_12580, n_12581, n_12582, n_12583, n_12584,
       n_12585;
  wire n_12586, n_12587, n_12588, n_12589, n_12590, n_12591, n_12592,
       n_12593;
  wire n_12594, n_12595, n_12596, n_12597, n_12598, n_12599, n_12600,
       n_12601;
  wire n_12602, n_12603, n_12604, n_12605, n_12606, n_12607, n_12608,
       n_12609;
  wire n_12610, n_12611, n_12612, n_12613, n_12614, n_12615, n_12616,
       n_12617;
  wire n_12618, n_12619, n_12620, n_12621, n_12622, n_12623, n_12624,
       n_12625;
  wire n_12626, n_12627, n_12628, n_12629, n_12630, n_12631, n_12632,
       n_12633;
  wire n_12634, n_12635, n_12636, n_12637, n_12638, n_12639, n_12640,
       n_12641;
  wire n_12642, n_12643, n_12644, n_12645, n_12646, n_12647, n_12648,
       n_12649;
  wire n_12650, n_12651, n_12652, n_12653, n_12654, n_12655, n_12656,
       n_12657;
  wire n_12658, n_12659, n_12660, n_12661, n_12662, n_12663, n_12664,
       n_12665;
  wire n_12666, n_12667, n_12668, n_12669, n_12670, n_12671, n_12672,
       n_12673;
  wire n_12674, n_12675, n_12676, n_12677, n_12678, n_12679, n_12680,
       n_12681;
  wire n_12682, n_12683, n_12684, n_12685, n_12686, n_12687, n_12688,
       n_12689;
  wire n_12690, n_12691, n_12692, n_12693, n_12694, n_12695, n_12696,
       n_12697;
  wire n_12698, n_12699, n_12700, n_12701, n_12702, n_12703, n_12704,
       n_12705;
  wire n_12706, n_12707, n_12708, n_12709, n_12710, n_12711, n_12712,
       n_12713;
  wire n_12714, n_12715, n_12716, n_12717, n_12718, n_12719, n_12720,
       n_12721;
  wire n_12722, n_12723, n_12724, n_12725, n_12726, n_12727, n_12728,
       n_12729;
  wire n_12730, n_12731, n_12732, n_12733, n_12734, n_12735, n_12736,
       n_12737;
  wire n_12738, n_12739, n_12740, n_12741, n_12742, n_12743, n_12744,
       n_12745;
  wire n_12746, n_12747, n_12748, n_12749, n_12750, n_12751, n_12752,
       n_12753;
  wire n_12754, n_12755, n_12756, n_12757, n_12758, n_12759, n_12760,
       n_12761;
  wire n_12762, n_12763, n_12764, n_12765, n_12766, n_12767, n_12768,
       n_12769;
  wire n_12770, n_12771, n_12772, n_12773, n_12774, n_12775, n_12776,
       n_12777;
  wire n_12778, n_12779, n_12780, n_12781, n_12782, n_12783, n_12784,
       n_12785;
  wire n_12786, n_12787, n_12788, n_12789, n_12790, n_12791, n_12792,
       n_12793;
  wire n_12794, n_12795, n_12796, n_12797, n_12798, n_12799, n_12800,
       n_12801;
  wire n_12802, n_12803, n_12804, n_12805, n_12806, n_12807, n_12808,
       n_12809;
  wire n_12810, n_12811, n_12812, n_12813, n_12814, n_12815, n_12816,
       n_12817;
  wire n_12818, n_12819, n_12820, n_12821, n_12822, n_12823, n_12824,
       n_12825;
  wire n_12826, n_12827, n_12828, n_12829, n_12830, n_12831, n_12832,
       n_12833;
  wire n_12834, n_12835, n_12836, n_12837, n_12838, n_12839, n_12840,
       n_12841;
  wire n_12842, n_12843, n_12844, n_12845, n_12846, n_12847, n_12848,
       n_12849;
  wire n_12850, n_12851, n_12852, n_12853, n_12854, n_12855, n_12856,
       n_12857;
  wire n_12858, n_12859, n_12860, n_12861, n_12862, n_12863, n_12864,
       n_12865;
  wire n_12866, n_12867, n_12868, n_12869, n_12870, n_12871, n_12872,
       n_12873;
  wire n_12874, n_12875, n_12876, n_12877, n_12878, n_12879, n_12880,
       n_12881;
  wire n_12882, n_12883, n_12884, n_12885, n_12886, n_12887, n_12888,
       n_12889;
  wire n_12890, n_12891, n_12892, n_12893, n_12894, n_12895, n_12896,
       n_12897;
  wire n_12898, n_12899, n_12900, n_12901, n_12902, n_12903, n_12904,
       n_12905;
  wire n_12906, n_12907, n_12908, n_12909, n_12910, n_12911, n_12912,
       n_12913;
  wire n_12914, n_12915, n_12916, n_12917, n_12918, n_12919, n_12920,
       n_12921;
  wire n_12922, n_12923, n_12924, n_12925, n_12926, n_12927, n_12928,
       n_12929;
  wire n_12930, n_12931, n_12932, n_12933, n_12934, n_12935, n_12936,
       n_12937;
  wire n_12938, n_12939, n_12940, n_12941, n_12942, n_12943, n_12944,
       n_12945;
  wire n_12946, n_12947, n_12948, n_12949, n_12950, n_12951, n_12952,
       n_12953;
  wire n_12954, n_12955, n_12956, n_12957, n_12958, n_12959, n_12960,
       n_12961;
  wire n_12962, n_12963, n_12964, n_12965, n_12966, n_12967, n_12968,
       n_12969;
  wire n_12970, n_12971, n_12972, n_12973, n_12974, n_12975, n_12976,
       n_12977;
  wire n_12978, n_12979, n_12980, n_12981, n_12982, n_12983, n_12984,
       n_12985;
  wire n_12986, n_12987, n_12988, n_12989, n_12990, n_12991, n_12992,
       n_12993;
  wire n_12994, n_12995, n_12996, n_12997, n_12998, n_12999, n_13000,
       n_13001;
  wire n_13002, n_13003, n_13004, n_13005, n_13006, n_13007, n_13008,
       n_13009;
  wire n_13010, n_13011, n_13012, n_13013, n_13014, n_13015, n_13016,
       n_13017;
  wire n_13018, n_13019, n_13020, n_13021, n_13022, n_13023, n_13024,
       n_13025;
  wire n_13026, n_13027, n_13028, n_13029, n_13030, n_13031, n_13032,
       n_13033;
  wire n_13034, n_13035, n_13036, n_13037, n_13038, n_13039, n_13040,
       n_13041;
  wire n_13042, n_13043, n_13044, n_13045, n_13046, n_13047, n_13048,
       n_13049;
  wire n_13050, n_13051, n_13052, n_13053, n_13054, n_13055, n_13056,
       n_13057;
  wire n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064,
       n_13065;
  wire n_13066, n_13067, n_13068, n_13069, n_13070, n_13071, n_13072,
       n_13073;
  wire n_13074, n_13075, n_13076, n_13077, n_13078, n_13079, n_13080,
       n_13081;
  wire n_13082, n_13083, n_13084, n_13085, n_13086, n_13087, n_13088,
       n_13089;
  wire n_13090, n_13091, n_13092, n_13093, n_13094, n_13095, n_13096,
       n_13097;
  wire n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104,
       n_13105;
  wire n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13112,
       n_13113;
  wire n_13114, n_13115, n_13116, n_13117, n_13118, n_13119, n_13120,
       n_13121;
  wire n_13122, n_13123, n_13124, n_13125, n_13126, n_13127, n_13128,
       n_13129;
  wire n_13130, n_13131, n_13132, n_13133, n_13134, n_13135, n_13136,
       n_13137;
  wire n_13138, n_13139, n_13140, n_13141, n_13142, n_13143, n_13144,
       n_13145;
  wire n_13146, n_13147, n_13148, n_13149, n_13150, n_13151, n_13152,
       n_13153;
  wire n_13154, n_13155, n_13156, n_13157, n_13158, n_13159, n_13160,
       n_13161;
  wire n_13162, n_13163, n_13164, n_13165, n_13166, n_13167, n_13168,
       n_13169;
  wire n_13170, n_13171, n_13172, n_13173, n_13174, n_13175, n_13176,
       n_13177;
  wire n_13178, n_13179, n_13180, n_13181, n_13182, n_13183, n_13184,
       n_13185;
  wire n_13186, n_13187, n_13188, n_13189, n_13190, n_13191, n_13192,
       n_13193;
  wire n_13194, n_13195, n_13196, n_13197, n_13198, n_13199, n_13200,
       n_13201;
  wire n_13202, n_13203, n_13204, n_13205, n_13206, n_13207, n_13208,
       n_13209;
  wire n_13210, n_13211, n_13212, n_13213, n_13214, n_13215, n_13216,
       n_13217;
  wire n_13218, n_13219, n_13220, n_13221, n_13222, n_13223, n_13224,
       n_13225;
  wire n_13226, n_13227, n_13228, n_13229, n_13230, n_13231, n_13232,
       n_13233;
  wire n_13234, n_13235, n_13236, n_13237, n_13238, n_13239, n_13240,
       n_13241;
  wire n_13242, n_13243, n_13244, n_13245, n_13246, n_13247, n_13248,
       n_13249;
  wire n_13250, n_13251, n_13252, n_13253, n_13254, n_13255, n_13256,
       n_13257;
  wire n_13258, n_13259, n_13260, n_13261, n_13262, n_13263, n_13264,
       n_13265;
  wire n_13266, n_13267, n_13268, n_13269, n_13270, n_13271, n_13272,
       n_13273;
  wire n_13274, n_13275, n_13276, n_13277, n_13278, n_13279, n_13280,
       n_13281;
  wire n_13282, n_13283, n_13284, n_13285, n_13286, n_13287, n_13288,
       n_13289;
  wire n_13290, n_13291, n_13292, n_13293, n_13294, n_13295, n_13296,
       n_13297;
  wire n_13298, n_13299, n_13300, n_13301, n_13302, n_13303, n_13304,
       n_13305;
  wire n_13306, n_13307, n_13308, n_13309, n_13310, n_13311, n_13312,
       n_13313;
  wire n_13314, n_13315, n_13316, n_13317, n_13318, n_13319, n_13320,
       n_13321;
  wire n_13322, n_13323, n_13324, n_13325, n_13326, n_13327, n_13328,
       n_13329;
  wire n_13330, n_13331, n_13332, n_13333, n_13334, n_13335, n_13336,
       n_13337;
  wire n_13338, n_13339, n_13340, n_13341, n_13342, n_13343, n_13344,
       n_13345;
  wire n_13346, n_13347, n_13348, n_13349, n_13350, n_13351, n_13352,
       n_13353;
  wire n_13354, n_13355, n_13356, n_13357, n_13358, n_13359, n_13360,
       n_13361;
  wire n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368,
       n_13369;
  wire n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376,
       n_13377;
  wire n_13378, n_13379, n_13380, n_13381, n_13382, n_13383, n_13384,
       n_13385;
  wire n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392,
       n_13393;
  wire n_13394, n_13395, n_13396, n_13397, n_13398, n_13399, n_13400,
       n_13401;
  wire n_13402, n_13403, n_13404, n_13405, n_13406, n_13407, n_13408,
       n_13409;
  wire n_13410, n_13411, n_13412, n_13413, n_13414, n_13415, n_13416,
       n_13417;
  wire n_13418, n_13419, n_13420, n_13421, n_13422, n_13423, n_13424,
       n_13425;
  wire n_13426, n_13427, n_13428, n_13429, n_13430, n_13431, n_13432,
       n_13433;
  wire n_13434, n_13435, n_13436, n_13437, n_13438, n_13439, n_13440,
       n_13441;
  wire n_13442, n_13443, n_13444, n_13445, n_13446, n_13447, n_13448,
       n_13449;
  wire n_13450, n_13451, n_13452, n_13453, n_13454, n_13455, n_13456,
       n_13457;
  wire n_13458, n_13459, n_13460, n_13461, n_13462, n_13463, n_13464,
       n_13465;
  wire n_13466, n_13467, n_13468, n_13469, n_13470, n_13471, n_13472,
       n_13473;
  wire n_13474, n_13475, n_13476, n_13477, n_13478, n_13479, n_13480,
       n_13481;
  wire n_13482, n_13483, n_13484, n_13485, n_13486, n_13487, n_13488,
       n_13489;
  wire n_13490, n_13491, n_13492, n_13493, n_13494, n_13495, n_13496,
       n_13497;
  wire n_13498, n_13499, n_13500, n_13501, n_13502, n_13503, n_13504,
       n_13505;
  wire n_13506, n_13507, n_13508, n_13509, n_13510, n_13511, n_13512,
       n_13513;
  wire n_13514, n_13515, n_13516, n_13517, n_13518, n_13519, n_13520,
       n_13521;
  wire n_13522, n_13523, n_13524, n_13525, n_13526, n_13527, n_13528,
       n_13529;
  wire n_13530, n_13531, n_13532, n_13533, n_13534, n_13535, n_13536,
       n_13537;
  wire n_13538, n_13539, n_13540, n_13541, n_13542, n_13543, n_13544,
       n_13545;
  wire n_13546, n_13547, n_13548, n_13549, n_13550, n_13551, n_13552,
       n_13553;
  wire n_13554, n_13555, n_13556, n_13557, n_13558, n_13559, n_13560,
       n_13561;
  wire n_13562, n_13563, n_13564, n_13565, n_13566, n_13567, n_13568,
       n_13569;
  wire n_13570, n_13571, n_13572, n_13573, n_13574, n_13575, n_13576,
       n_13577;
  wire n_13578, n_13579, n_13580, n_13581, n_13582, n_13583, n_13584,
       n_13585;
  wire n_13586, n_13587, n_13588, n_13589, n_13590, n_13591, n_13592,
       n_13593;
  wire n_13594, n_13595, n_13596, n_13597, n_13598, n_13599, n_13600,
       n_13601;
  wire n_13602, n_13603, n_13604, n_13605, n_13606, n_13607, n_13608,
       n_13609;
  wire n_13610, n_13611, n_13612, n_13613, n_13614, n_13615, n_13616,
       n_13617;
  wire n_13618, n_13619, n_13620, n_13621, n_13622, n_13623, n_13624,
       n_13625;
  wire n_13626, n_13627, n_13628, n_13629, n_13630, n_13631, n_13632,
       n_13633;
  wire n_13634, n_13635, n_13636, n_13637, n_13638, n_13639, n_13640,
       n_13641;
  wire n_13642, n_13643, n_13644, n_13645, n_13646, n_13647, n_13648,
       n_13649;
  wire n_13650, n_13651, n_13652, n_13653, n_13654, n_13655, n_13656,
       n_13657;
  wire n_13658, n_13659, n_13660, n_13661, n_13662, n_13663, n_13664,
       n_13665;
  wire n_13666, n_13667, n_13668, n_13669, n_13670, n_13671, n_13672,
       n_13673;
  wire n_13674, n_13675, n_13676, n_13677, n_13678, n_13679, n_13680,
       n_13681;
  wire n_13682, n_13683, n_13684, n_13685, n_13686, n_13687, n_13688,
       n_13689;
  wire n_13690, n_13691, n_13692, n_13693, n_13694, n_13695, n_13696,
       n_13697;
  wire n_13698, n_13699, n_13700, n_13701, n_13702, n_13703, n_13704,
       n_13705;
  wire n_13706, n_13707, n_13708, n_13709, n_13710, n_13711, n_13712,
       n_13713;
  wire n_13714, n_13715, n_13716, n_13717, n_13718, n_13719, n_13720,
       n_13721;
  wire n_13722, n_13723, n_13724, n_13725, n_13726, n_13727, n_13728,
       n_13729;
  wire n_13730, n_13731, n_13732, n_13733, n_13734, n_13735, n_13736,
       n_13737;
  wire n_13738, n_13739, n_13740, n_13741, n_13742, n_13743, n_13744,
       n_13745;
  wire n_13746, n_13747, n_13748, n_13749, n_13750, n_13751, n_13752,
       n_13753;
  wire n_13754, n_13755, n_13756, n_13757, n_13758, n_13759, n_13760,
       n_13761;
  wire n_13762, n_13763, n_13764, n_13765, n_13766, n_13767, n_13768,
       n_13769;
  wire n_13770, n_13771, n_13772, n_13773, n_13774, n_13775, n_13776,
       n_13777;
  wire n_13778, n_13779, n_13780, n_13781, n_13782, n_13783, n_13784,
       n_13785;
  wire n_13786, n_13787, n_13788, n_13789, n_13790, n_13791, n_13792,
       n_13793;
  wire n_13794, n_13795, n_13796, n_13797, n_13798, n_13799, n_13800,
       n_13801;
  wire n_13802, n_13803, n_13804, n_13805, n_13806, n_13807, n_13808,
       n_13809;
  wire n_13810, n_13811, n_13812, n_13813, n_13814, n_13815, n_13816,
       n_13817;
  wire n_13818, n_13819, n_13820, n_13821, n_13822, n_13823, n_13824,
       n_13825;
  wire n_13826, n_13827, n_13828, n_13829, n_13830, n_13831, n_13832,
       n_13833;
  wire n_13834, n_13835, n_13836, n_13837, n_13838, n_13839, n_13840,
       n_13841;
  wire n_13842, n_13843, n_13844, n_13845, n_13846, n_13847, n_13848,
       n_13849;
  wire n_13850, n_13851, n_13852, n_13853, n_13854, n_13855, n_13856,
       n_13857;
  wire n_13858, n_13859, n_13860, n_13861, n_13862, n_13863, n_13864,
       n_13865;
  wire n_13866, n_13867, n_13868, n_13869, n_13870, n_13871, n_13872,
       n_13873;
  wire n_13874, n_13875, n_13876, n_13877, n_13878, n_13879, n_13880,
       n_13881;
  wire n_13882, n_13883, n_13884, n_13885, n_13886, n_13887, n_13888,
       n_13889;
  wire n_13890, n_13891, n_13892, n_13893, n_13894, n_13895, n_13896,
       n_13897;
  wire n_13898, n_13899, n_13900, n_13901, n_13902, n_13903, n_13904,
       n_13905;
  wire n_13906, n_13907, n_13908, n_13909, n_13910, n_13911, n_13912,
       n_13913;
  wire n_13914, n_13915, n_13916, n_13917, n_13918, n_13919, n_13920,
       n_13921;
  wire n_13922, n_13923, n_13924, n_13925, n_13926, n_13927, n_13928,
       n_13929;
  wire n_13930, n_13931, n_13932, n_13933, n_13934, n_13935, n_13936,
       n_13937;
  wire n_13938, n_13939, n_13940, n_13941, n_13942, n_13943, n_13944,
       n_13945;
  wire n_13946, n_13947, n_13948, n_13949, n_13950, n_13951, n_13952,
       n_13953;
  wire n_13954, n_13955, n_13956, n_13957, n_13958, n_13959, n_13960,
       n_13961;
  wire n_13962, n_13963, n_13964, n_13965, n_13966, n_13967, n_13968,
       n_13969;
  wire n_13970, n_13971, n_13972, n_13973, n_13974, n_13975, n_13976,
       n_13977;
  wire n_13978, n_13979, n_13980, n_13981, n_13982, n_13983, n_13984,
       n_13985;
  wire n_13986, n_13987, n_13988, n_13989, n_13990, n_13991, n_13992,
       n_13993;
  wire n_13994, n_13995, n_13996, n_13997, n_13998, n_13999, n_14000,
       n_14001;
  wire n_14002, n_14003, n_14004, n_14005, n_14006, n_14007, n_14008,
       n_14009;
  wire n_14010, n_14011, n_14012, n_14013, n_14014, n_14015, n_14016,
       n_14017;
  wire n_14018, n_14019, n_14020, n_14021, n_14022, n_14023, n_14024,
       n_14025;
  wire n_14026, n_14027, n_14028, n_14029, n_14030, n_14031, n_14032,
       n_14033;
  wire n_14034, n_14035, n_14036, n_14037, n_14038, n_14039, n_14040,
       n_14041;
  wire n_14042, n_14043, n_14044, n_14045, n_14046, n_14047, n_14048,
       n_14049;
  wire n_14050, n_14051, n_14052, n_14053, n_14054, n_14055, n_14056,
       n_14057;
  wire n_14058, n_14059, n_14060, n_14061, n_14062, n_14063, n_14064,
       n_14065;
  wire n_14066, n_14067, n_14068, n_14069, n_14070, n_14071, n_14072,
       n_14073;
  wire n_14074, n_14075, n_14076, n_14077, n_14078, n_14079, n_14080,
       n_14081;
  wire n_14082, n_14083, n_14084, n_14085, n_14086, n_14087, n_14088,
       n_14089;
  wire n_14090, n_14091, n_14092, n_14093, n_14094, n_14095, n_14096,
       n_14097;
  wire n_14098, n_14099, n_14100, n_14101, n_14102, n_14103, n_14104,
       n_14105;
  wire n_14106, n_14107, n_14108, n_14109, n_14110, n_14111, n_14112,
       n_14113;
  wire n_14114, n_14115, n_14116, n_14117, n_14118, n_14119, n_14120,
       n_14121;
  wire n_14122, n_14123, n_14124, n_14125, n_14126, n_14127, n_14128,
       n_14129;
  wire n_14130, n_14131, n_14132, n_14133, n_14134, n_14135, n_14136,
       n_14137;
  wire n_14138, n_14139, n_14140, n_14141, n_14142, n_14143, n_14144,
       n_14145;
  wire n_14146, n_14147, n_14148, n_14149, n_14150, n_14151, n_14152,
       n_14153;
  wire n_14154, n_14155, n_14156, n_14157, n_14158, n_14159, n_14160,
       n_14161;
  wire n_14162, n_14163, n_14164, n_14165, n_14166, n_14167, n_14168,
       n_14169;
  wire n_14170, n_14171, n_14172, n_14173, n_14174, n_14175, n_14176,
       n_14177;
  wire n_14178, n_14179, n_14180, n_14181, n_14182, n_14183, n_14184,
       n_14185;
  wire n_14186, n_14187, n_14188, n_14189, n_14190, n_14191, n_14192,
       n_14193;
  wire n_14194, n_14195, n_14196, n_14197, n_14198, n_14199, n_14200,
       n_14201;
  wire n_14202, n_14203, n_14204, n_14205, n_14206, n_14207, n_14208,
       n_14209;
  wire n_14210, n_14211, n_14212, n_14213, n_14214, n_14215, n_14216,
       n_14217;
  wire n_14218, n_14219, n_14220, n_14221, n_14222, n_14223, n_14224,
       n_14225;
  wire n_14226, n_14227, n_14228, n_14229, n_14230, n_14231, n_14232,
       n_14233;
  wire n_14234, n_14235, n_14236, n_14237, n_14238, n_14239, n_14240,
       n_14241;
  wire n_14242, n_14243, n_14244, n_14245, n_14246, n_14247, n_14248,
       n_14249;
  wire n_14250, n_14251, n_14252, n_14253, n_14254, n_14255, n_14256,
       n_14257;
  wire n_14258, n_14259, n_14260, n_14261, n_14262, n_14263, n_14264,
       n_14265;
  wire n_14266, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272,
       n_14273;
  wire n_14274, n_14275, n_14276, n_14277, n_14278, n_14279, n_14280,
       n_14281;
  wire n_14282, n_14283, n_14284, n_14285, n_14286, n_14287, n_14288,
       n_14289;
  wire n_14290, n_14291, n_14292, n_14293, n_14294, n_14295, n_14296,
       n_14297;
  wire n_14298, n_14299, n_14300, n_14301, n_14302, n_14303, n_14304,
       n_14305;
  wire n_14306, n_14307, n_14308, n_14309, n_14310, n_14311, n_14312,
       n_14313;
  wire n_14314, n_14315, n_14316, n_14317, n_14318, n_14319, n_14320,
       n_14321;
  wire n_14322, n_14323, n_14324, n_14325, n_14326, n_14327, n_14328,
       n_14329;
  wire n_14330, n_14331, n_14332, n_14333, n_14334, n_14335, n_14336,
       n_14337;
  wire n_14338, n_14339, n_14340, n_14341, n_14342, n_14343, n_14344,
       n_14345;
  wire n_14346, n_14347, n_14348, n_14349, n_14350, n_14351, n_14352,
       n_14353;
  wire n_14354, n_14355, n_14356, n_14357, n_14358, n_14359, n_14360,
       n_14361;
  wire n_14362, n_14363, n_14364, n_14365, n_14366, n_14367, n_14368,
       n_14369;
  wire n_14370, n_14371, n_14372, n_14373, n_14374, n_14375, n_14376,
       n_14377;
  wire n_14378, n_14379, n_14380, n_14381, n_14382, n_14383, n_14384,
       n_14385;
  wire n_14386, n_14387, n_14388, n_14389, n_14390, n_14391, n_14392,
       n_14393;
  wire n_14394, n_14395, n_14396, n_14397, n_14398, n_14399, n_14400,
       n_14401;
  wire n_14402, n_14403, n_14404, n_14405, n_14406, n_14407, n_14408,
       n_14409;
  wire n_14410, n_14411, n_14412, n_14413, n_14414, n_14415, n_14416,
       n_14417;
  wire n_14418, n_14419, n_14420, n_14421, n_14422, n_14423, n_14424,
       n_14425;
  wire n_14426, n_14427, n_14428, n_14429, n_14430, n_14431, n_14432,
       n_14433;
  wire n_14434, n_14435, n_14436, n_14437, n_14438, n_14439, n_14440,
       n_14441;
  wire n_14442, n_14443, n_14444, n_14445, n_14446, n_14447, n_14448,
       n_14449;
  wire n_14450, n_14451, n_14452, n_14453, n_14454, n_14455, n_14456,
       n_14457;
  wire n_14458, n_14459, n_14460, n_14461, n_14462, n_14463, n_14464,
       n_14465;
  wire n_14466, n_14467, n_14468, n_14469, n_14470, n_14471, n_14472,
       n_14473;
  wire n_14474, n_14475, n_14476, n_14477, n_14478, n_14479, n_14480,
       n_14481;
  wire n_14482, n_14483, n_14484, n_14485, n_14486, n_14487, n_14488,
       n_14489;
  wire n_14490, n_14491, n_14492, n_14493, n_14494, n_14495, n_14496,
       n_14497;
  wire n_14498, n_14499, n_14500, n_14501, n_14502, n_14503, n_14504,
       n_14505;
  wire n_14506, n_14507, n_14508, n_14509, n_14510, n_14511, n_14512,
       n_14513;
  wire n_14514, n_14515, n_14516, n_14517, n_14518, n_14519, n_14520,
       n_14521;
  wire n_14522, n_14523, n_14524, n_14525, n_14526, n_14527, n_14528,
       n_14529;
  wire n_14530, n_14531, n_14532, n_14533, n_14534, n_14535, n_14536,
       n_14537;
  wire n_14538, n_14539, n_14540, n_14541, n_14542, n_14543, n_14544,
       n_14545;
  wire n_14546, n_14547, n_14548, n_14549, n_14550, n_14551, n_14552,
       n_14553;
  wire n_14554, n_14555, n_14556, n_14557, n_14558, n_14559, n_14560,
       n_14561;
  wire n_14562, n_14563, n_14564, n_14565, n_14566, n_14567, n_14568,
       n_14569;
  wire n_14570, n_14571, n_14572, n_14573, n_14574, n_14575, n_14576,
       n_14577;
  wire n_14578, n_14579, n_14580, n_14581, n_14582, n_14583, n_14584,
       n_14585;
  wire n_14586, n_14587, n_14588, n_14589, n_14590, n_14591, n_14592,
       n_14593;
  wire n_14594, n_14595, n_14596, n_14597, n_14598, n_14599, n_14600,
       n_14601;
  wire n_14602, n_14603, n_14604, n_14605, n_14606, n_14607, n_14608,
       n_14609;
  wire n_14610, n_14611, n_14612, n_14613, n_14614, n_14615, n_14616,
       n_14617;
  wire n_14618, n_14619, n_14620, n_14621, n_14622, n_14623, n_14624,
       n_14625;
  wire n_14626, n_14627, n_14628, n_14629, n_14630, n_14631, n_14632,
       n_14633;
  wire n_14634, n_14635, n_14636, n_14637, n_14638, n_14639, n_14640,
       n_14641;
  wire n_14642, n_14643, n_14644, n_14645, n_14646, n_14647, n_14648,
       n_14649;
  wire n_14650, n_14651, n_14652, n_14653, n_14654, n_14655, n_14656,
       n_14657;
  wire n_14658, n_14659, n_14660, n_14661, n_14662, n_14663, n_14664,
       n_14665;
  wire n_14666, n_14667, n_14668, n_14669, n_14670, n_14671, n_14672,
       n_14673;
  wire n_14674, n_14675, n_14676, n_14677, n_14678, n_14679, n_14680,
       n_14681;
  wire n_14682, n_14683, n_14684, n_14685, n_14686, n_14687, n_14688,
       n_14689;
  wire n_14690, n_14691, n_14692, n_14693, n_14694, n_14695, n_14696,
       n_14697;
  wire n_14698, n_14699, n_14700, n_14701, n_14702, n_14703, n_14704,
       n_14705;
  wire n_14706, n_14707, n_14708, n_14709, n_14710, n_14711, n_14712,
       n_14713;
  wire n_14714, n_14715, n_14716, n_14717, n_14718, n_14719, n_14720,
       n_14721;
  wire n_14722, n_14723, n_14724, n_14725, n_14726, n_14727, n_14728,
       n_14729;
  wire n_14730, n_14731, n_14732, n_14733, n_14734, n_14735, n_14736,
       n_14737;
  wire n_14738, n_14739, n_14740, n_14741, n_14742, n_14743, n_14744,
       n_14745;
  wire n_14746, n_14747, n_14748, n_14749, n_14750, n_14751, n_14752,
       n_14753;
  wire n_14754, n_14755, n_14756, n_14757, n_14758, n_14759, n_14760,
       n_14761;
  wire n_14762, n_14763, n_14764, n_14765, n_14766, n_14767, n_14768,
       n_14769;
  wire n_14770, n_14771, n_14772, n_14773, n_14774, n_14775, n_14776,
       n_14777;
  wire n_14778, n_14779, n_14780, n_14781, n_14782, n_14783, n_14784,
       n_14785;
  wire n_14786, n_14787, n_14788, n_14789, n_14790, n_14791, n_14792,
       n_14793;
  wire n_14794, n_14795, n_14796, n_14797, n_14798, n_14799, n_14800,
       n_14801;
  wire n_14802, n_14803, n_14804, n_14805, n_14806, n_14807, n_14808,
       n_14809;
  wire n_14810, n_14811, n_14812, n_14813, n_14814, n_14815, n_14816,
       n_14817;
  wire n_14818, n_14819, n_14820, n_14821, n_14822, n_14823, n_14824,
       n_14825;
  wire n_14826, n_14827, n_14828, n_14829, n_14830, n_14831, n_14832,
       n_14833;
  wire n_14834, n_14835, n_14836, n_14837, n_14838, n_14839, n_14840,
       n_14841;
  wire n_14842, n_14843, n_14844, n_14845, n_14846, n_14847, n_14848,
       n_14849;
  wire n_14850, n_14851, n_14852, n_14853, n_14854, n_14855, n_14856,
       n_14857;
  wire n_14858, n_14859, n_14860, n_14861, n_14862, n_14863, n_14864,
       n_14865;
  wire n_14866, n_14867, n_14868, n_14869, n_14870, n_14871, n_14872,
       n_14873;
  wire n_14874, n_14875, n_14876, n_14877, n_14878, n_14879, n_14880,
       n_14881;
  wire n_14882, n_14883, n_14884, n_14885, n_14886, n_14887, n_14888,
       n_14889;
  wire n_14890, n_14891, n_14892, n_14893, n_14894, n_14895, n_14896,
       n_14897;
  wire n_14898, n_14899, n_14900, n_14901, n_14902, n_14903, n_14904,
       n_14905;
  wire n_14906, n_14907, n_14908, n_14909, n_14910, n_14911, n_14912,
       n_14913;
  wire n_14914, n_14915, n_14916, n_14917, n_14918, n_14919, n_14920,
       n_14921;
  wire n_14922, n_14923, n_14924, n_14925, n_14926, n_14927, n_14928,
       n_14929;
  wire n_14930, n_14931, n_14932, n_14933, n_14934, n_14935, n_14936,
       n_14937;
  wire n_14938, n_14939, n_14940, n_14941, n_14942, n_14943, n_14944,
       n_14945;
  wire n_14946, n_14947, n_14948, n_14949, n_14950, n_14951, n_14952,
       n_14953;
  wire n_14954, n_14955, n_14956, n_14957, n_14958, n_14959, n_14960,
       n_14961;
  wire n_14962, n_14963, n_14964, n_14965, n_14966, n_14967, n_14968,
       n_14969;
  wire n_14970, n_14971, n_14972, n_14973, n_14974, n_14975, n_14976,
       n_14977;
  wire n_14978, n_14979, n_14980, n_14981, n_14982, n_14983, n_14984,
       n_14985;
  wire n_14986, n_14987, n_14988, n_14989, n_14990, n_14991, n_14992,
       n_14993;
  wire n_14994, n_14995, n_14996, n_14997, n_14998, n_14999, n_15000,
       n_15001;
  wire n_15002, n_15003, n_15004, n_15005, n_15006, n_15007, n_15008,
       n_15009;
  wire n_15010, n_15011, n_15012, n_15013, n_15014, n_15015, n_15016,
       n_15017;
  wire n_15018, n_15019, n_15020, n_15021, n_15022, n_15023, n_15024,
       n_15025;
  wire n_15026, n_15027, n_15028, n_15029, n_15030, n_15031, n_15032,
       n_15033;
  wire n_15034, n_15035, n_15036, n_15037, n_15038, n_15039, n_15040,
       n_15041;
  wire n_15042, n_15043, n_15044, n_15045, n_15046, n_15047, n_15048,
       n_15049;
  wire n_15050, n_15051, n_15052, n_15053, n_15054, n_15055, n_15056,
       n_15057;
  wire n_15058, n_15059, n_15060, n_15061, n_15062, n_15063, n_15064,
       n_15065;
  wire n_15066, n_15067, n_15068, n_15069, n_15070, n_15071, n_15072,
       n_15073;
  wire n_15074, n_15075, n_15076, n_15077, n_15078, n_15079, n_15080,
       n_15081;
  wire n_15082, n_15083, n_15084, n_15085, n_15086, n_15087, n_15088,
       n_15089;
  wire n_15090, n_15091, n_15092, n_15093, n_15094, n_15095, n_15096,
       n_15097;
  wire n_15098, n_15099, n_15100, n_15101, n_15102, n_15103, n_15104,
       n_15105;
  wire n_15106, n_15107, n_15108, n_15109, n_15110, n_15111, n_15112,
       n_15113;
  wire n_15114, n_15115, n_15116, n_15117, n_15118, n_15119, n_15120,
       n_15121;
  wire n_15122, n_15123, n_15124, n_15125, n_15126, n_15127, n_15128,
       n_15129;
  wire n_15130, n_15131, n_15132, n_15133, n_15134, n_15135, n_15136,
       n_15137;
  wire n_15138, n_15139, n_15140, n_15141, n_15142, n_15143, n_15144,
       n_15145;
  wire n_15146, n_15147, n_15148, n_15149, n_15150, n_15151, n_15152,
       n_15153;
  wire n_15154, n_15155, n_15156, n_15157, n_15158, n_15159, n_15160,
       n_15161;
  wire n_15162, n_15163, n_15164, n_15165, n_15166, n_15167, n_15168,
       n_15169;
  wire n_15170, n_15171, n_15172, n_15173, n_15174, n_15175, n_15176,
       n_15177;
  wire n_15178, n_15179, n_15180, n_15181, n_15182, n_15183, n_15184,
       n_15185;
  wire n_15186, n_15187, n_15188, n_15189, n_15190, n_15191, n_15192,
       n_15193;
  wire n_15194, n_15195, n_15196, n_15197, n_15198, n_15199, n_15200,
       n_15201;
  wire n_15202, n_15203, n_15204, n_15205, n_15206, n_15207, n_15208,
       n_15209;
  wire n_15210, n_15211, n_15212, n_15213, n_15214, n_15215, n_15216,
       n_15217;
  wire n_15218, n_15219, n_15220, n_15221, n_15222, n_15223, n_15224,
       n_15225;
  wire n_15226, n_15227, n_15228, n_15229, n_15230, n_15231, n_15232,
       n_15233;
  wire n_15234, n_15235, n_15236, n_15237, n_15238, n_15239, n_15240,
       n_15241;
  wire n_15242, n_15243, n_15244, n_15245, n_15246, n_15247, n_15248,
       n_15249;
  wire n_15250, n_15251, n_15252, n_15253, n_15254, n_15255, n_15256,
       n_15257;
  wire n_15258, n_15259, n_15260, n_15261, n_15262, n_15263, n_15264,
       n_15265;
  wire n_15266, n_15267, n_15268, n_15269, n_15270, n_15271, n_15272,
       n_15273;
  wire n_15274, n_15275, n_15276, n_15277, n_15278, n_15279, n_15280,
       n_15281;
  wire n_15282, n_15283, n_15284, n_15285, n_15286, n_15287, n_15288,
       n_15289;
  wire n_15290, n_15291, n_15292, n_15293, n_15294, n_15295, n_15296,
       n_15297;
  wire n_15298, n_15299, n_15300, n_15301, n_15302, n_15303, n_15304,
       n_15305;
  wire n_15306, n_15307, n_15308, n_15309, n_15310, n_15311, n_15312,
       n_15313;
  wire n_15314, n_15315, n_15316, n_15317, n_15318, n_15319, n_15320,
       n_15321;
  wire n_15322, n_15323, n_15324, n_15325, n_15326, n_15327, n_15328,
       n_15329;
  wire n_15330, n_15331, n_15332, n_15333, n_15334, n_15335, n_15336,
       n_15337;
  wire n_15338, n_15339, n_15340, n_15341, n_15342, n_15343, n_15344,
       n_15345;
  wire n_15346, n_15347, n_15348, n_15349, n_15350, n_15351, n_15352,
       n_15353;
  wire n_15354, n_15355, n_15356, n_15357, n_15358, n_15359, n_15360,
       n_15361;
  wire n_15362, n_15363, n_15364, n_15365, n_15366, n_15367, n_15368,
       n_15369;
  wire n_15370, n_15371, n_15372, n_15373, n_15374, n_15375, n_15376,
       n_15377;
  wire n_15378, n_15379, n_15380, n_15381, n_15382, n_15383, n_15384,
       n_15385;
  wire n_15386, n_15387, n_15388, n_15389, n_15390, n_15391, n_15392,
       n_15393;
  wire n_15394, n_15395, n_15396, n_15397, n_15398, n_15399, n_15400,
       n_15401;
  wire n_15402, n_15403, n_15404, n_15405, n_15406, n_15407, n_15408,
       n_15409;
  wire n_15410, n_15411, n_15412, n_15413, n_15414, n_15415, n_15416,
       n_15417;
  wire n_15418, n_15419, n_15420, n_15421, n_15422, n_15423, n_15424,
       n_15425;
  wire n_15426, n_15427, n_15428, n_15429, n_15430, n_15431, n_15432,
       n_15433;
  wire n_15434, n_15435, n_15436, n_15437, n_15438, n_15439, n_15440,
       n_15441;
  wire n_15442, n_15443, n_15444, n_15445, n_15446, n_15447, n_15448,
       n_15449;
  wire n_15450, n_15451, n_15452, n_15453, n_15454, n_15455, n_15456,
       n_15457;
  wire n_15458, n_15459, n_15460, n_15461, n_15462, n_15463, n_15464,
       n_15465;
  wire n_15466, n_15467, n_15468, n_15469, n_15470, n_15471, n_15472,
       n_15473;
  wire n_15474, n_15475, n_15476, n_15477, n_15478, n_15479, n_15480,
       n_15481;
  wire n_15482, n_15483, n_15484, n_15485, n_15486, n_15487, n_15488,
       n_15489;
  wire n_15490, n_15491, n_15492, n_15493, n_15494, n_15495, n_15496,
       n_15497;
  wire n_15498, n_15499, n_15500, n_15501, n_15502, n_15503, n_15504,
       n_15505;
  wire n_15506, n_15507, n_15508, n_15509, n_15510, n_15511, n_15512,
       n_15513;
  wire n_15514, n_15515, n_15516, n_15517, n_15518, n_15519, n_15520,
       n_15521;
  wire n_15522, n_15523, n_15524, n_15525, n_15526, n_15527, n_15528,
       n_15529;
  wire n_15530, n_15531, n_15532, n_15533, n_15534, n_15535, n_15536,
       n_15537;
  wire n_15538, n_15539, n_15540, n_15541, n_15542, n_15543, n_15544,
       n_15545;
  wire n_15546, n_15547, n_15548, n_15549, n_15550, n_15551, n_15552,
       n_15553;
  wire n_15554, n_15555, n_15556, n_15557, n_15558, n_15559, n_15560,
       n_15561;
  wire n_15562, n_15563, n_15564, n_15565, n_15566, n_15567, n_15568,
       n_15569;
  wire n_15570, n_15571, n_15572, n_15573, n_15574, n_15575, n_15576,
       n_15577;
  wire n_15578, n_15579, n_15580, n_15581, n_15582, n_15583, n_15584,
       n_15585;
  wire n_15586, n_15587, n_15588, n_15589, n_15590, n_15591, n_15592,
       n_15593;
  wire n_15594, n_15595, n_15596, n_15597, n_15598, n_15599, n_15600,
       n_15601;
  wire n_15602, n_15603, n_15604, n_15605, n_15606, n_15607, n_15608,
       n_15609;
  wire n_15610, n_15611, n_15612, n_15613, n_15614, n_15615, n_15616,
       n_15617;
  wire n_15618, n_15619, n_15620, n_15621, n_15622, n_15623, n_15624,
       n_15625;
  wire n_15626, n_15627, n_15628, n_15629, n_15630, n_15631, n_15632,
       n_15633;
  wire n_15634, n_15635, n_15636, n_15637, n_15638, n_15639, n_15640,
       n_15641;
  wire n_15642, n_15643, n_15644, n_15645, n_15646, n_15647, n_15648,
       n_15649;
  wire n_15650, n_15651, n_15652, n_15653, n_15654, n_15655, n_15656,
       n_15657;
  wire n_15658, n_15659, n_15660, n_15661, n_15662, n_15663, n_15664,
       n_15665;
  wire n_15666, n_15667, n_15668, n_15669, n_15670, n_15671, n_15672,
       n_15673;
  wire n_15674, n_15675, n_15676, n_15677, n_15678, n_15679, n_15680,
       n_15681;
  wire n_15682, n_15683, n_15684, n_15685, n_15686, n_15687, n_15688,
       n_15689;
  wire n_15690, n_15691, n_15692, n_15693, n_15694, n_15695, n_15696,
       n_15697;
  wire n_15698, n_15699, n_15700, n_15701, n_15702, n_15703, n_15704,
       n_15705;
  wire n_15706, n_15707, n_15708, n_15709, n_15710, n_15711, n_15712,
       n_15713;
  wire n_15714, n_15715, n_15716, n_15717, n_15718, n_15719, n_15720,
       n_15721;
  wire n_15722, n_15723, n_15724, n_15725, n_15726, n_15727, n_15728,
       n_15729;
  wire n_15730, n_15731, n_15732, n_15733, n_15734, n_15735, n_15736,
       n_15737;
  wire n_15738, n_15739, n_15740, n_15741, n_15742, n_15743, n_15744,
       n_15745;
  wire n_15746, n_15747, n_15748, n_15749, n_15750, n_15751, n_15752,
       n_15753;
  wire n_15754, n_15755, n_15756, n_15757, n_15758, n_15759, n_15760,
       n_15761;
  wire n_15762, n_15763, n_15764, n_15765, n_15766, n_15767, n_15768,
       n_15769;
  wire n_15770, n_15771, n_15772, n_15773, n_15774, n_15775, n_15776,
       n_15777;
  wire n_15778, n_15779, n_15780, n_15781, n_15782, n_15783, n_15784,
       n_15785;
  wire n_15786, n_15787, n_15788, n_15789, n_15790, n_15791, n_15792,
       n_15793;
  wire n_15794, n_15795, n_15796, n_15797, n_15798, n_15799, n_15800,
       n_15801;
  wire n_15802, n_15803, n_15804, n_15805, n_15806, n_15807, n_15808,
       n_15809;
  wire n_15810, n_15811, n_15812, n_15813, n_15814, n_15815, n_15816,
       n_15817;
  wire n_15818, n_15819, n_15820, n_15821, n_15822, n_15823, n_15824,
       n_15825;
  wire n_15826, n_15827, n_15828, n_15829, n_15830, n_15831, n_15832,
       n_15833;
  wire n_15834, n_15835, n_15836, n_15837, n_15838, n_15839, n_15840,
       n_15841;
  wire n_15842, n_15843, n_15844, n_15845, n_15846, n_15847, n_15848,
       n_15849;
  wire n_15850, n_15851, n_15852, n_15853, n_15854, n_15855, n_15856,
       n_15857;
  wire n_15858, n_15859, n_15860, n_15861, n_15862, n_15863, n_15864,
       n_15865;
  wire n_15866, n_15867, n_15868, n_15869, n_15870, n_15871, n_15872,
       n_15873;
  wire n_15874, n_15875, n_15876, n_15877, n_15878, n_15879, n_15880,
       n_15881;
  wire n_15882, n_15883, n_15884, n_15885, n_15886, n_15887, n_15888,
       n_15889;
  wire n_15890, n_15891, n_15892, n_15893, n_15894, n_15895, n_15896,
       n_15897;
  wire n_15898, n_15899, n_15900, n_15901, n_15902, n_15903, n_15904,
       n_15905;
  wire n_15906, n_15907, n_15908, n_15909, n_15910, n_15911, n_15912,
       n_15913;
  wire n_15914, n_15915, n_15916, n_15917, n_15918, n_15919, n_15920,
       n_15921;
  wire n_15922, n_15923, n_15924, n_15925, n_15926, n_15927, n_15928,
       n_15929;
  wire n_15930, n_15931, n_15932, n_15933, n_15934, n_15935, n_15936,
       n_15937;
  wire n_15938, n_15939, n_15940, n_15941, n_15942, n_15943, n_15944,
       n_15945;
  wire n_15946, n_15947, n_15948, n_15949, n_15950, n_15951, n_15952,
       n_15953;
  wire n_15954, n_15955, n_15956, n_15957, n_15958, n_15959, n_15960,
       n_15961;
  wire n_15962, n_15963, n_15964, n_15965, n_15966, n_15967, n_15968,
       n_15969;
  wire n_15970, n_15971, n_15972, n_15973, n_15974, n_15975, n_15976,
       n_15977;
  wire n_15978, n_15979, n_15980, n_15981, n_15982, n_15983, n_15984,
       n_15985;
  wire n_15986, n_15987, n_15988, n_15989, n_15990, n_15991, n_15992,
       n_15993;
  wire n_15994, n_15995, n_15996, n_15997, n_15998, n_15999, n_16000,
       n_16001;
  wire n_16002, n_16003, n_16004, n_16005, n_16006, n_16007, n_16008,
       n_16009;
  wire n_16010, n_16011, n_16012, n_16013, n_16014, n_16015, n_16016,
       n_16017;
  wire n_16018, n_16019, n_16020, n_16021, n_16022, n_16023, n_16024,
       n_16025;
  wire n_16026, n_16027, n_16028, n_16029, n_16030, n_16031, n_16032,
       n_16033;
  wire n_16034, n_16035, n_16036, n_16037, n_16038, n_16039, n_16040,
       n_16041;
  wire n_16042, n_16043, n_16044, n_16045, n_16046, n_16047, n_16048,
       n_16049;
  wire n_16050, n_16051, n_16052, n_16053, n_16054, n_16055, n_16056,
       n_16057;
  wire n_16058, n_16059, n_16060, n_16061, n_16062, n_16063, n_16064,
       n_16065;
  wire n_16066, n_16067, n_16068, n_16069, n_16070, n_16071, n_16072,
       n_16073;
  wire n_16074, n_16075, n_16076, n_16077, n_16078, n_16079, n_16080,
       n_16081;
  wire n_16082, n_16083, n_16084, n_16085, n_16086, n_16087, n_16088,
       n_16089;
  wire n_16090, n_16091, n_16092, n_16093, n_16094, n_16095, n_16096,
       n_16097;
  wire n_16098, n_16099, n_16100, n_16101, n_16102, n_16103, n_16104,
       n_16105;
  wire n_16106, n_16107, n_16108, n_16109, n_16110, n_16111, n_16112,
       n_16113;
  wire n_16114, n_16115, n_16116, n_16117, n_16118, n_16119, n_16120,
       n_16121;
  wire n_16122, n_16123, n_16124, n_16125, n_16126, n_16127, n_16128,
       n_16129;
  wire n_16130, n_16131, n_16132, n_16133, n_16134, n_16135, n_16136,
       n_16137;
  wire n_16138, n_16139, n_16140, n_16141, n_16142, n_16143, n_16144,
       n_16145;
  wire n_16146, n_16147, n_16148, n_16149, n_16150, n_16151, n_16152,
       n_16153;
  wire n_16154, n_16155, n_16156, n_16157, n_16158, n_16159, n_16160,
       n_16161;
  wire n_16162, n_16163, n_16164, n_16165, n_16166, n_16167, n_16168,
       n_16169;
  wire n_16170, n_16171, n_16172, n_16173, n_16174, n_16175, n_16176,
       n_16177;
  wire n_16178, n_16179, n_16180, n_16181, n_16182, n_16183, n_16184,
       n_16185;
  wire n_16186, n_16187, n_16188, n_16189, n_16190, n_16191, n_16192,
       n_16193;
  wire n_16194, n_16195, n_16196, n_16197, n_16198, n_16199, n_16200,
       n_16201;
  wire n_16202, n_16203, n_16204, n_16205, n_16206, n_16207, n_16208,
       n_16209;
  wire n_16210, n_16211, n_16212, n_16213, n_16214, n_16215, n_16216,
       n_16217;
  wire n_16218, n_16219, n_16220, n_16221, n_16222, n_16223, n_16224,
       n_16225;
  wire n_16226, n_16227, n_16228, n_16229, n_16230, n_16231, n_16232,
       n_16233;
  wire n_16234, n_16235, n_16236, n_16237, n_16238, n_16239, n_16240,
       n_16241;
  wire n_16242, n_16243, n_16244, n_16245, n_16246, n_16247, n_16248,
       n_16249;
  wire n_16250, n_16251, n_16252, n_16253, n_16254, n_16255, n_16256,
       n_16257;
  wire n_16258, n_16259, n_16260, n_16261, n_16262, n_16263, n_16264,
       n_16265;
  wire n_16266, n_16267, n_16268, n_16269, n_16270, n_16271, n_16272,
       n_16273;
  wire n_16274, n_16275, n_16276, n_16277, n_16278, n_16279, n_16280,
       n_16281;
  wire n_16282, n_16283, n_16284, n_16285, n_16286, n_16287, n_16288,
       n_16289;
  wire n_16290, n_16291, n_16292, n_16293, n_16294, n_16295, n_16296,
       n_16297;
  wire n_16298, n_16299, n_16300, n_16301, n_16302, n_16303, n_16304,
       n_16305;
  wire n_16306, n_16307, n_16308, n_16309, n_16310, n_16311, n_16312,
       n_16313;
  wire n_16314, n_16315, n_16316, n_16317, n_16318, n_16319, n_16320,
       n_16321;
  wire n_16322, n_16323, n_16324, n_16325, n_16326, n_16327, n_16328,
       n_16329;
  wire n_16330, n_16331, n_16332, n_16333, n_16334, n_16335, n_16336,
       n_16337;
  wire n_16338, n_16339, n_16340, n_16341, n_16342, n_16343, n_16344,
       n_16345;
  wire n_16346, n_16347, n_16348, n_16349, n_16350, n_16351, n_16352,
       n_16353;
  wire n_16354, n_16355, n_16356, n_16357, n_16358, n_16359, n_16360,
       n_16361;
  wire n_16362, n_16363, n_16364, n_16365, n_16366, n_16367, n_16368,
       n_16369;
  wire n_16370, n_16371, n_16372, n_16373, n_16374, n_16375, n_16376,
       n_16377;
  wire n_16378, n_16379, n_16380, n_16381, n_16382, n_16383, n_16384,
       n_16385;
  wire n_16386, n_16387, n_16388, n_16389, n_16390, n_16391, n_16392,
       n_16393;
  wire n_16394, n_16395, n_16396, n_16397, n_16398, n_16399, n_16400,
       n_16401;
  wire n_16402, n_16403, n_16404, n_16405, n_16406, n_16407, n_16408,
       n_16409;
  wire n_16410, n_16411, n_16412, n_16413, n_16414, n_16415, n_16416,
       n_16417;
  wire n_16418, n_16419, n_16420, n_16421, n_16422, n_16423, n_16424,
       n_16425;
  wire n_16426, n_16427, n_16428, n_16429, n_16430, n_16431, n_16432,
       n_16433;
  wire n_16434, n_16435, n_16436, n_16437, n_16438, n_16439, n_16440,
       n_16441;
  wire n_16442, n_16443, n_16444, n_16445, n_16446, n_16447, n_16448,
       n_16449;
  wire n_16450, n_16451, n_16452, n_16453, n_16454, n_16455, n_16456,
       n_16457;
  wire n_16458, n_16459, n_16460, n_16461, n_16462, n_16463, n_16464,
       n_16465;
  wire n_16466, n_16467, n_16468, n_16469, n_16470, n_16471, n_16472,
       n_16473;
  wire n_16474, n_16475, n_16476, n_16477, n_16478, n_16479, n_16480,
       n_16481;
  wire n_16482, n_16483, n_16484, n_16485, n_16486, n_16487, n_16488,
       n_16489;
  wire n_16490, n_16491, n_16492, n_16493, n_16494, n_16495, n_16496,
       n_16497;
  wire n_16498, n_16499, n_16500, n_16501, n_16502, n_16503, n_16504,
       n_16505;
  wire n_16506, n_16507, n_16508, n_16509, n_16510, n_16511, n_16512,
       n_16513;
  wire n_16514, n_16515, n_16516, n_16517, n_16518, n_16519, n_16520,
       n_16521;
  wire n_16522, n_16523, n_16524, n_16525, n_16526, n_16527, n_16528,
       n_16529;
  wire n_16530, n_16531, n_16532, n_16533, n_16534, n_16535, n_16536,
       n_16537;
  wire n_16538, n_16539, n_16540, n_16541, n_16542, n_16543, n_16544,
       n_16545;
  wire n_16546, n_16547, n_16548, n_16549, n_16550, n_16551, n_16552,
       n_16553;
  wire n_16554, n_16555, n_16556, n_16557, n_16558, n_16559, n_16560,
       n_16561;
  wire n_16562, n_16563, n_16564, n_16565, n_16566, n_16567, n_16568,
       n_16569;
  wire n_16570, n_16571, n_16572, n_16573, n_16574, n_16575, n_16576,
       n_16577;
  wire n_16578, n_16579, n_16580, n_16581, n_16582, n_16583, n_16584,
       n_16585;
  wire n_16586, n_16587, n_16588, n_16589, n_16590, n_16591, n_16592,
       n_16593;
  wire n_16594, n_16595, n_16596, n_16597, n_16598, n_16599, n_16600,
       n_16601;
  wire n_16602, n_16603, n_16604, n_16605, n_16606, n_16607, n_16608,
       n_16609;
  wire n_16610, n_16611, n_16612, n_16613, n_16614, n_16615, n_16616,
       n_16617;
  wire n_16618, n_16619, n_16620, n_16621, n_16622, n_16623, n_16624,
       n_16625;
  wire n_16626, n_16627, n_16628, n_16629, n_16630, n_16631, n_16632,
       n_16633;
  wire n_16634, n_16635, n_16636, n_16637, n_16638, n_16639, n_16640,
       n_16641;
  wire n_16642, n_16643, n_16644, n_16645, n_16646, n_16647, n_16648,
       n_16649;
  wire n_16650, n_16651, n_16652, n_16653, n_16654, n_16655, n_16656,
       n_16657;
  wire n_16658, n_16659, n_16660, n_16661, n_16662, n_16663, n_16664,
       n_16665;
  wire n_16666, n_16667, n_16668, n_16669, n_16670, n_16671, n_16672,
       n_16673;
  wire n_16674, n_16675, n_16676, n_16677, n_16678, n_16679, n_16680,
       n_16681;
  wire n_16682, n_16683, n_16684, n_16685, n_16686, n_16687, n_16688,
       n_16689;
  wire n_16690, n_16691, n_16692, n_16693, n_16694, n_16695, n_16696,
       n_16697;
  wire n_16698, n_16699, n_16700, n_16701, n_16702, n_16703, n_16704,
       n_16705;
  wire n_16706, n_16707, n_16708, n_16709, n_16710, n_16711, n_16712,
       n_16713;
  wire n_16714, n_16715, n_16716, n_16717, n_16718, n_16719, n_16720,
       n_16721;
  wire n_16722, n_16723, n_16724, n_16725, n_16726, n_16727, n_16728,
       n_16729;
  wire n_16730, n_16731, n_16732, n_16733, n_16734, n_16735, n_16736,
       n_16737;
  wire n_16738, n_16739, n_16740, n_16741, n_16742, n_16743, n_16744,
       n_16745;
  wire n_16746, n_16747, n_16748, n_16749, n_16750, n_16751, n_16752,
       n_16753;
  wire n_16754, n_16755, n_16756, n_16757, n_16758, n_16759, n_16760,
       n_16761;
  wire n_16762, n_16763, n_16764, n_16765, n_16766, n_16767, n_16768,
       n_16769;
  wire n_16770, n_16771, n_16772, n_16773, n_16774, n_16775, n_16776,
       n_16777;
  wire n_16778, n_16779, n_16780, n_16781, n_16782, n_16783, n_16784,
       n_16785;
  wire n_16786, n_16787, n_16788, n_16789, n_16790, n_16791, n_16792,
       n_16793;
  wire n_16794, n_16795, n_16796, n_16797, n_16798, n_16799, n_16800,
       n_16801;
  wire n_16802, n_16803, n_16804, n_16805, n_16806, n_16807, n_16808,
       n_16809;
  wire n_16810, n_16811, n_16812, n_16813, n_16814, n_16815, n_16816,
       n_16817;
  wire n_16818, n_16819, n_16820, n_16821, n_16822, n_16823, n_16824,
       n_16825;
  wire n_16826, n_16827, n_16828, n_16829, n_16830, n_16831, n_16832,
       n_16833;
  wire n_16834, n_16835, n_16836, n_16837, n_16838, n_16839, n_16840,
       n_16841;
  wire n_16842, n_16843, n_16844, n_16845, n_16846, n_16847, n_16848,
       n_16849;
  wire n_16850, n_16851, n_16852, n_16853, n_16854, n_16855, n_16856,
       n_16857;
  wire n_16858, n_16859, n_16860, n_16861, n_16862, n_16863, n_16864,
       n_16865;
  wire n_16866, n_16867, n_16868, n_16869, n_16870, n_16871, n_16872,
       n_16873;
  wire n_16874, n_16875, n_16876, n_16877, n_16878, n_16879, n_16880,
       n_16881;
  wire n_16882, n_16883, n_16884, n_16885, n_16886, n_16887, n_16888,
       n_16889;
  wire n_16890, n_16891, n_16892, n_16893, n_16894, n_16895, n_16896,
       n_16897;
  wire n_16898, n_16899, n_16900, n_16901, n_16902, n_16903, n_16904,
       n_16905;
  wire n_16906, n_16907, n_16908, n_16909, n_16910, n_16911, n_16912,
       n_16913;
  wire n_16914, n_16915, n_16916, n_16917, n_16918, n_16919, n_16920,
       n_16921;
  wire n_16922, n_16923, n_16924, n_16925, n_16926, n_16927, n_16928,
       n_16929;
  wire n_16930, n_16931, n_16932, n_16933, n_16934, n_16935, n_16936,
       n_16937;
  wire n_16938, n_16939, n_16940, n_16941, n_16942, n_16943, n_16944,
       n_16945;
  wire n_16946, n_16947, n_16948, n_16949, n_16950, n_16951, n_16952,
       n_16953;
  wire n_16954, n_16955, n_16956, n_16957, n_16958, n_16959, n_16960,
       n_16961;
  wire n_16962, n_16963, n_16964, n_16965, n_16966, n_16967, n_16968,
       n_16969;
  wire n_16970, n_16971, n_16972, n_16973, n_16974, n_16975, n_16976,
       n_16977;
  wire n_16978, n_16979, n_16980, n_16981, n_16982, n_16983, n_16984,
       n_16985;
  wire n_16986, n_16987, n_16988, n_16989, n_16990, n_16991, n_16992,
       n_16993;
  wire n_16994, n_16995, n_16996, n_16997, n_16998, n_16999, n_17000,
       n_17001;
  wire n_17002, n_17003, n_17004, n_17005, n_17006, n_17007, n_17008,
       n_17009;
  wire n_17010, n_17011, n_17012, n_17013, n_17014, n_17015, n_17016,
       n_17017;
  wire n_17018, n_17019, n_17020, n_17021, n_17022, n_17023, n_17024,
       n_17025;
  wire n_17026, n_17027, n_17028, n_17029, n_17030, n_17031, n_17032,
       n_17033;
  wire n_17034, n_17035, n_17036, n_17037, n_17038, n_17039, n_17040,
       n_17041;
  wire n_17042, n_17043, n_17044, n_17045, n_17046, n_17047, n_17048,
       n_17049;
  wire n_17050, n_17051, n_17052, n_17053, n_17054, n_17055, n_17056,
       n_17057;
  wire n_17058, n_17059, n_17060, n_17061, n_17062, n_17063, n_17064,
       n_17065;
  wire n_17066, n_17067, n_17068, n_17069, n_17070, n_17071, n_17072,
       n_17073;
  assign \asquared[1]  = 1'b0;
  assign \asquared[0]  = \a[0] ;
  and g1 (n194, \a[0] , \a[1] );
  not g2 (n_4, n194);
  and g3 (\asquared[2] , \a[1] , n_4);
  and g4 (n196, \a[0] , \a[2] );
  and g5 (n197, n194, n196);
  not g6 (n_6, n196);
  and g7 (n198, n_4, n_6);
  not g8 (n_7, n197);
  not g9 (n_8, n198);
  and g10 (\asquared[3] , n_7, n_8);
  and g11 (n200, \a[1] , \a[2] );
  not g12 (n_9, n200);
  and g13 (n201, \a[2] , n_9);
  and g14 (n202, \a[0] , \a[3] );
  not g15 (n_11, n201);
  not g16 (n_12, n202);
  and g17 (n203, n_11, n_12);
  and g18 (n204, n201, n202);
  not g19 (n_13, n203);
  not g20 (n_14, n204);
  and g21 (n205, n_13, n_14);
  not g22 (n_15, n205);
  and g23 (n206, n197, n_15);
  and g24 (n207, n_7, n205);
  or g25 (\asquared[4] , n206, n207);
  and g26 (n209, \a[3] , \a[4] );
  and g27 (n210, n194, n209);
  and g28 (n211, \a[1] , \a[3] );
  and g29 (n212, \a[0] , \a[4] );
  not g30 (n_17, n211);
  not g31 (n_18, n212);
  and g32 (n213, n_17, n_18);
  not g33 (n_19, n210);
  not g34 (n_20, n213);
  and g35 (n214, n_19, n_20);
  not g36 (n_21, n214);
  and g37 (n215, n_9, n_21);
  and g38 (n216, n200, n214);
  not g39 (n_22, n215);
  not g40 (n_23, n216);
  and g41 (n217, n_22, n_23);
  and g42 (n218, \a[2] , \a[3] );
  and g43 (n219, \a[0] , n218);
  not g44 (n_24, n217);
  not g45 (n_25, n219);
  and g46 (n220, n_24, n_25);
  and g47 (n221, n217, n219);
  not g48 (n_26, n220);
  not g49 (n_27, n221);
  and g50 (\asquared[5] , n_26, n_27);
  and g51 (n223, \a[1] , \a[4] );
  and g52 (n224, \a[0] , \a[5] );
  not g53 (n_29, n223);
  not g54 (n_30, n224);
  and g55 (n225, n_29, n_30);
  and g56 (n226, \a[4] , \a[5] );
  and g57 (n227, n194, n226);
  not g58 (n_31, n225);
  not g59 (n_32, n227);
  and g60 (n228, n_31, n_32);
  and g61 (n229, n210, n228);
  not g62 (n_33, n229);
  and g63 (n230, n_32, n_33);
  and g64 (n231, n_31, n230);
  and g65 (n232, n210, n_33);
  not g66 (n_34, n231);
  not g67 (n_35, n232);
  and g68 (n233, n_34, n_35);
  not g69 (n_36, n218);
  and g70 (n234, \a[3] , n_36);
  not g71 (n_37, n234);
  and g72 (n235, n233, n_37);
  not g73 (n_38, n233);
  and g74 (n236, n_38, n234);
  not g75 (n_39, n235);
  not g76 (n_40, n236);
  and g77 (n237, n_39, n_40);
  and g78 (n238, n_22, n219);
  not g79 (n_41, n238);
  and g80 (n239, n_23, n_41);
  not g81 (n_42, n237);
  and g82 (n240, n_42, n239);
  not g83 (n_43, n239);
  and g84 (n241, n237, n_43);
  not g85 (n_44, n240);
  not g86 (n_45, n241);
  and g87 (\asquared[6] , n_44, n_45);
  and g88 (n243, n_39, n_43);
  not g89 (n_46, n243);
  and g90 (n244, n_40, n_46);
  and g91 (n245, \a[6] , n219);
  not g92 (n_48, n245);
  and g93 (n246, \a[0] , n_48);
  and g94 (n247, \a[6] , n246);
  and g95 (n248, n218, n_48);
  not g96 (n_49, n247);
  not g97 (n_50, n248);
  and g98 (n249, n_49, n_50);
  and g99 (n250, n200, n226);
  and g100 (n251, \a[1] , \a[5] );
  and g101 (n252, \a[2] , \a[4] );
  not g102 (n_51, n251);
  not g103 (n_52, n252);
  and g104 (n253, n_51, n_52);
  not g105 (n_53, n250);
  not g106 (n_54, n253);
  and g107 (n254, n_53, n_54);
  not g108 (n_55, n254);
  and g109 (n255, n249, n_55);
  not g110 (n_56, n249);
  and g111 (n256, n_56, n254);
  not g112 (n_57, n255);
  not g113 (n_58, n256);
  and g114 (n257, n_57, n_58);
  not g115 (n_59, n257);
  and g116 (n258, n230, n_59);
  not g117 (n_60, n230);
  and g118 (n259, n_60, n257);
  not g119 (n_61, n258);
  not g120 (n_62, n259);
  and g121 (n260, n_61, n_62);
  not g122 (n_63, n260);
  and g123 (n261, n244, n_63);
  not g124 (n_64, n244);
  and g125 (n262, n_64, n_61);
  and g126 (n263, n_62, n262);
  not g127 (n_65, n261);
  not g128 (n_66, n263);
  and g129 (\asquared[7] , n_65, n_66);
  and g130 (n265, n218, n226);
  and g131 (n266, \a[0] , \a[7] );
  and g132 (n267, n209, n266);
  and g133 (n268, \a[5] , \a[7] );
  and g134 (n269, n196, n268);
  not g135 (n_68, n267);
  not g136 (n_69, n269);
  and g137 (n270, n_68, n_69);
  not g138 (n_70, n265);
  not g139 (n_71, n270);
  and g140 (n271, n_70, n_71);
  not g141 (n_72, n271);
  and g142 (n272, n_70, n_72);
  and g143 (n273, \a[2] , \a[5] );
  not g144 (n_73, n209);
  not g145 (n_74, n273);
  and g146 (n274, n_73, n_74);
  not g147 (n_75, n274);
  and g148 (n275, n272, n_75);
  and g149 (n276, n266, n_72);
  not g150 (n_76, n275);
  not g151 (n_77, n276);
  and g152 (n277, n_76, n_77);
  and g153 (n278, n_48, n_58);
  and g154 (n279, \a[1] , \a[6] );
  not g155 (n_78, n279);
  and g156 (n280, n250, n_78);
  not g157 (n_79, n280);
  and g158 (n281, n250, n_79);
  not g159 (n_80, \a[4] );
  and g160 (n282, n_80, n_78);
  and g161 (n283, \a[4] , n279);
  not g162 (n_81, n283);
  and g163 (n284, n_79, n_81);
  not g164 (n_82, n282);
  and g165 (n285, n_82, n284);
  not g166 (n_83, n281);
  not g167 (n_84, n285);
  and g168 (n286, n_83, n_84);
  not g169 (n_85, n278);
  not g170 (n_86, n286);
  and g171 (n287, n_85, n_86);
  and g172 (n288, n278, n_84);
  and g173 (n289, n_83, n288);
  not g174 (n_87, n287);
  not g175 (n_88, n289);
  and g176 (n290, n_87, n_88);
  not g177 (n_89, n290);
  and g178 (n291, n277, n_89);
  not g179 (n_90, n277);
  and g180 (n292, n_90, n290);
  not g181 (n_91, n291);
  not g182 (n_92, n292);
  and g183 (n293, n_91, n_92);
  not g184 (n_93, n262);
  and g185 (n294, n_62, n_93);
  not g186 (n_94, n293);
  and g187 (n295, n_94, n294);
  not g188 (n_95, n294);
  and g189 (n296, n293, n_95);
  not g190 (n_96, n295);
  not g191 (n_97, n296);
  and g192 (\asquared[8] , n_96, n_97);
  and g193 (n298, n_79, n_87);
  and g194 (n299, \a[1] , \a[7] );
  and g195 (n300, \a[3] , \a[5] );
  and g196 (n301, n299, n300);
  not g197 (n_98, n301);
  and g198 (n302, n299, n_98);
  and g199 (n303, n300, n_98);
  not g200 (n_99, n302);
  not g201 (n_100, n303);
  and g202 (n304, n_99, n_100);
  not g203 (n_101, n272);
  not g204 (n_102, n304);
  and g205 (n305, n_101, n_102);
  not g206 (n_103, n305);
  and g207 (n306, n_101, n_103);
  and g208 (n307, n_102, n_103);
  not g209 (n_104, n306);
  not g210 (n_105, n307);
  and g211 (n308, n_104, n_105);
  and g212 (n309, \a[0] , \a[8] );
  and g213 (n310, \a[2] , \a[6] );
  not g214 (n_107, n309);
  not g215 (n_108, n310);
  and g216 (n311, n_107, n_108);
  and g217 (n312, \a[6] , \a[8] );
  and g218 (n313, n196, n312);
  not g219 (n_109, n311);
  not g220 (n_110, n313);
  and g221 (n314, n_109, n_110);
  and g222 (n315, n283, n314);
  not g223 (n_111, n315);
  and g224 (n316, n_110, n_111);
  and g225 (n317, n_109, n316);
  and g226 (n318, n283, n_111);
  not g227 (n_112, n317);
  not g228 (n_113, n318);
  and g229 (n319, n_112, n_113);
  not g230 (n_114, n308);
  not g231 (n_115, n319);
  and g232 (n320, n_114, n_115);
  and g233 (n321, n308, n319);
  not g234 (n_116, n320);
  not g235 (n_117, n321);
  and g236 (n322, n_116, n_117);
  not g237 (n_118, n322);
  and g238 (n323, n298, n_118);
  not g239 (n_119, n298);
  and g240 (n324, n_119, n322);
  not g241 (n_120, n323);
  not g242 (n_121, n324);
  and g243 (n325, n_120, n_121);
  and g244 (n326, n_91, n_95);
  not g245 (n_122, n326);
  and g246 (n327, n_92, n_122);
  not g247 (n_123, n325);
  and g248 (n328, n_123, n327);
  not g249 (n_124, n327);
  and g250 (n329, n325, n_124);
  not g251 (n_125, n328);
  not g252 (n_126, n329);
  and g253 (\asquared[9] , n_125, n_126);
  and g254 (n331, n_103, n_116);
  and g255 (n332, \a[5] , \a[6] );
  and g256 (n333, n209, n332);
  and g257 (n334, n252, n268);
  and g258 (n335, \a[6] , \a[7] );
  and g259 (n336, n218, n335);
  not g260 (n_127, n334);
  not g261 (n_128, n336);
  and g262 (n337, n_127, n_128);
  not g263 (n_129, n333);
  not g264 (n_130, n337);
  and g265 (n338, n_129, n_130);
  not g266 (n_131, n338);
  and g267 (n339, n_129, n_131);
  and g268 (n340, \a[3] , \a[6] );
  not g269 (n_132, n226);
  not g270 (n_133, n340);
  and g271 (n341, n_132, n_133);
  not g272 (n_134, n341);
  and g273 (n342, n339, n_134);
  and g274 (n343, \a[2] , \a[7] );
  and g275 (n344, n_131, n343);
  not g276 (n_135, n342);
  not g277 (n_136, n344);
  and g278 (n345, n_135, n_136);
  not g279 (n_137, n316);
  not g280 (n_138, n345);
  and g281 (n346, n_137, n_138);
  not g282 (n_139, n346);
  and g283 (n347, n_137, n_139);
  and g284 (n348, n_138, n_139);
  not g285 (n_140, n347);
  not g286 (n_141, n348);
  and g287 (n349, n_140, n_141);
  and g288 (n350, \a[0] , \a[9] );
  not g289 (n_143, n350);
  and g290 (n351, n301, n_143);
  and g291 (n352, n_98, n350);
  not g292 (n_144, n351);
  not g293 (n_145, n352);
  and g294 (n353, n_144, n_145);
  and g295 (n354, \a[5] , \a[8] );
  and g296 (n355, \a[1] , n354);
  not g297 (n_146, n355);
  and g298 (n356, \a[5] , n_146);
  and g299 (n357, \a[1] , n_146);
  and g300 (n358, \a[8] , n357);
  not g301 (n_147, n356);
  not g302 (n_148, n358);
  and g303 (n359, n_147, n_148);
  not g304 (n_149, n353);
  not g305 (n_150, n359);
  and g306 (n360, n_149, n_150);
  and g307 (n361, n353, n359);
  not g308 (n_151, n360);
  not g309 (n_152, n361);
  and g310 (n362, n_151, n_152);
  not g311 (n_153, n349);
  and g312 (n363, n_153, n362);
  not g313 (n_154, n362);
  and g314 (n364, n_141, n_154);
  and g315 (n365, n_140, n364);
  not g316 (n_155, n363);
  not g317 (n_156, n365);
  and g318 (n366, n_155, n_156);
  not g319 (n_157, n331);
  and g320 (n367, n_157, n366);
  not g321 (n_158, n366);
  and g322 (n368, n331, n_158);
  not g323 (n_159, n367);
  not g324 (n_160, n368);
  and g325 (n369, n_159, n_160);
  and g326 (n370, n_120, n_124);
  not g327 (n_161, n370);
  and g328 (n371, n_121, n_161);
  not g329 (n_162, n369);
  and g330 (n372, n_162, n371);
  not g331 (n_163, n371);
  and g332 (n373, n369, n_163);
  not g333 (n_164, n372);
  not g334 (n_165, n373);
  and g335 (\asquared[10] , n_164, n_165);
  and g336 (n375, n_160, n_163);
  not g337 (n_166, n375);
  and g338 (n376, n_159, n_166);
  and g339 (n377, n_139, n_155);
  and g340 (n378, \a[8] , \a[10] );
  and g341 (n379, n196, n378);
  and g342 (n380, \a[7] , \a[8] );
  and g343 (n381, n218, n380);
  not g344 (n_168, n379);
  not g345 (n_169, n381);
  and g346 (n382, n_168, n_169);
  and g347 (n383, \a[0] , \a[10] );
  and g348 (n384, \a[3] , \a[7] );
  and g349 (n385, n383, n384);
  not g350 (n_170, n382);
  not g351 (n_171, n385);
  and g352 (n386, n_170, n_171);
  not g353 (n_172, n386);
  and g354 (n387, \a[2] , n_172);
  and g355 (n388, \a[8] , n387);
  and g356 (n389, n_171, n_172);
  not g357 (n_173, n383);
  not g358 (n_174, n384);
  and g359 (n390, n_173, n_174);
  not g360 (n_175, n390);
  and g361 (n391, n389, n_175);
  not g362 (n_176, n388);
  not g363 (n_177, n391);
  and g364 (n392, n_176, n_177);
  and g365 (n393, n301, n350);
  not g366 (n_178, n393);
  and g367 (n394, n_151, n_178);
  not g368 (n_179, n392);
  and g369 (n395, n_179, n394);
  not g370 (n_180, n394);
  and g371 (n396, n392, n_180);
  not g372 (n_181, n395);
  not g373 (n_182, n396);
  and g374 (n397, n_181, n_182);
  and g375 (n398, \a[9] , n283);
  and g376 (n399, \a[1] , \a[9] );
  and g377 (n400, \a[4] , \a[6] );
  not g378 (n_183, n399);
  not g379 (n_184, n400);
  and g380 (n401, n_183, n_184);
  not g381 (n_185, n398);
  not g382 (n_186, n401);
  and g383 (n402, n_185, n_186);
  and g384 (n403, n355, n402);
  not g385 (n_187, n403);
  and g386 (n404, n355, n_187);
  and g387 (n405, n402, n_187);
  not g388 (n_188, n404);
  not g389 (n_189, n405);
  and g390 (n406, n_188, n_189);
  not g391 (n_190, n339);
  not g392 (n_191, n406);
  and g393 (n407, n_190, n_191);
  and g394 (n408, n339, n_189);
  and g395 (n409, n_188, n408);
  not g396 (n_192, n407);
  not g397 (n_193, n409);
  and g398 (n410, n_192, n_193);
  not g399 (n_194, n397);
  and g400 (n411, n_194, n410);
  not g401 (n_195, n410);
  and g402 (n412, n397, n_195);
  not g403 (n_196, n411);
  not g404 (n_197, n412);
  and g405 (n413, n_196, n_197);
  not g406 (n_198, n413);
  and g407 (n414, n377, n_198);
  not g408 (n_199, n377);
  and g409 (n415, n_199, n413);
  not g410 (n_200, n414);
  not g411 (n_201, n415);
  and g412 (n416, n_200, n_201);
  not g413 (n_202, n416);
  and g414 (n417, n376, n_202);
  not g415 (n_203, n376);
  and g416 (n418, n_203, n_200);
  and g417 (n419, n_201, n418);
  not g418 (n_204, n417);
  not g419 (n_205, n419);
  and g420 (\asquared[11] , n_204, n_205);
  and g421 (n421, n_179, n_180);
  not g422 (n_206, n421);
  and g423 (n422, n_196, n_206);
  and g424 (n423, \a[10] , n279);
  not g425 (n_207, n423);
  and g426 (n424, \a[6] , n_207);
  and g427 (n425, \a[1] , n_207);
  and g428 (n426, \a[10] , n425);
  not g429 (n_208, n424);
  not g430 (n_209, n426);
  and g431 (n427, n_208, n_209);
  not g432 (n_210, n389);
  not g433 (n_211, n427);
  and g434 (n428, n_210, n_211);
  not g435 (n_212, n428);
  and g436 (n429, n_210, n_212);
  and g437 (n430, n_211, n_212);
  not g438 (n_213, n429);
  not g439 (n_214, n430);
  and g440 (n431, n_213, n_214);
  and g441 (n432, \a[8] , \a[9] );
  and g442 (n433, n218, n432);
  and g443 (n434, \a[2] , \a[9] );
  and g444 (n435, \a[3] , \a[8] );
  not g445 (n_215, n434);
  not g446 (n_216, n435);
  and g447 (n436, n_215, n_216);
  not g448 (n_217, n433);
  not g449 (n_218, n436);
  and g450 (n437, n_217, n_218);
  and g451 (n438, n398, n437);
  not g452 (n_219, n438);
  and g453 (n439, n398, n_219);
  and g454 (n440, n_217, n_219);
  and g455 (n441, n_218, n440);
  not g456 (n_220, n439);
  not g457 (n_221, n441);
  and g458 (n442, n_220, n_221);
  not g459 (n_222, n431);
  not g460 (n_223, n442);
  and g461 (n443, n_222, n_223);
  not g462 (n_224, n443);
  and g463 (n444, n_222, n_224);
  and g464 (n445, n_223, n_224);
  not g465 (n_225, n444);
  not g466 (n_226, n445);
  and g467 (n446, n_225, n_226);
  and g468 (n447, n_187, n_192);
  and g469 (n448, n226, n335);
  and g470 (n449, \a[0] , \a[11] );
  and g471 (n450, \a[4] , \a[7] );
  not g472 (n_228, n332);
  not g473 (n_229, n450);
  and g474 (n451, n_228, n_229);
  not g475 (n_230, n448);
  not g476 (n_231, n451);
  and g477 (n452, n_230, n_231);
  and g478 (n453, n449, n452);
  not g479 (n_232, n453);
  and g480 (n454, n_230, n_232);
  and g481 (n455, n_231, n454);
  and g482 (n456, n449, n_232);
  not g483 (n_233, n455);
  not g484 (n_234, n456);
  and g485 (n457, n_233, n_234);
  not g486 (n_235, n447);
  not g487 (n_236, n457);
  and g488 (n458, n_235, n_236);
  not g489 (n_237, n458);
  and g490 (n459, n_235, n_237);
  and g491 (n460, n_236, n_237);
  not g492 (n_238, n459);
  not g493 (n_239, n460);
  and g494 (n461, n_238, n_239);
  not g495 (n_240, n446);
  not g496 (n_241, n461);
  and g497 (n462, n_240, n_241);
  and g498 (n463, n446, n_239);
  and g499 (n464, n_238, n463);
  not g500 (n_242, n462);
  not g501 (n_243, n464);
  and g502 (n465, n_242, n_243);
  not g503 (n_244, n465);
  and g504 (n466, n422, n_244);
  not g505 (n_245, n422);
  and g506 (n467, n_245, n465);
  not g507 (n_246, n466);
  not g508 (n_247, n467);
  and g509 (n468, n_246, n_247);
  not g510 (n_248, n418);
  and g511 (n469, n_201, n_248);
  not g512 (n_249, n468);
  and g513 (n470, n_249, n469);
  not g514 (n_250, n469);
  and g515 (n471, n468, n_250);
  not g516 (n_251, n470);
  not g517 (n_252, n471);
  and g518 (\asquared[12] , n_251, n_252);
  and g519 (n473, n_246, n_250);
  not g520 (n_253, n473);
  and g521 (n474, n_247, n_253);
  and g522 (n475, n_237, n_242);
  and g523 (n476, n440, n454);
  not g524 (n_254, n440);
  not g525 (n_255, n454);
  and g526 (n477, n_254, n_255);
  not g527 (n_256, n476);
  not g528 (n_257, n477);
  and g529 (n478, n_256, n_257);
  and g530 (n479, \a[3] , \a[9] );
  and g531 (n480, \a[10] , \a[12] );
  and g532 (n481, n196, n480);
  and g533 (n482, \a[0] , \a[12] );
  and g534 (n483, n479, n482);
  and g535 (n484, \a[9] , \a[10] );
  and g536 (n485, n218, n484);
  not g537 (n_259, n483);
  not g538 (n_260, n485);
  and g539 (n486, n_259, n_260);
  not g540 (n_261, n481);
  not g541 (n_262, n486);
  and g542 (n487, n_261, n_262);
  not g543 (n_263, n487);
  and g544 (n488, n479, n_263);
  and g545 (n489, n_261, n_263);
  and g546 (n490, \a[2] , \a[10] );
  not g547 (n_264, n482);
  not g548 (n_265, n490);
  and g549 (n491, n_264, n_265);
  not g550 (n_266, n491);
  and g551 (n492, n489, n_266);
  not g552 (n_267, n488);
  not g553 (n_268, n492);
  and g554 (n493, n_267, n_268);
  not g555 (n_269, n493);
  and g556 (n494, n478, n_269);
  not g557 (n_270, n494);
  and g558 (n495, n478, n_270);
  and g559 (n496, n_269, n_270);
  not g560 (n_271, n495);
  not g561 (n_272, n496);
  and g562 (n497, n_271, n_272);
  and g563 (n498, n_212, n_224);
  and g564 (n499, \a[4] , \a[8] );
  not g565 (n_273, n499);
  and g566 (n500, n_207, n_273);
  and g567 (n501, n423, n499);
  and g568 (n502, \a[5] , \a[11] );
  and g569 (n503, n299, n502);
  and g570 (n504, \a[1] , \a[11] );
  not g571 (n_274, n268);
  not g572 (n_275, n504);
  and g573 (n505, n_274, n_275);
  not g574 (n_276, n503);
  not g575 (n_277, n505);
  and g576 (n506, n_276, n_277);
  not g577 (n_278, n501);
  and g578 (n507, n_278, n506);
  not g579 (n_279, n500);
  and g580 (n508, n_279, n507);
  not g581 (n_280, n508);
  and g582 (n509, n_278, n_280);
  and g583 (n510, n_279, n509);
  and g584 (n511, n506, n_280);
  not g585 (n_281, n510);
  not g586 (n_282, n511);
  and g587 (n512, n_281, n_282);
  not g588 (n_283, n498);
  not g589 (n_284, n512);
  and g590 (n513, n_283, n_284);
  and g591 (n514, n498, n512);
  not g592 (n_285, n513);
  not g593 (n_286, n514);
  and g594 (n515, n_285, n_286);
  not g595 (n_287, n497);
  and g596 (n516, n_287, n515);
  not g597 (n_288, n515);
  and g598 (n517, n497, n_288);
  not g599 (n_289, n516);
  not g600 (n_290, n517);
  and g601 (n518, n_289, n_290);
  not g602 (n_291, n518);
  and g603 (n519, n475, n_291);
  not g604 (n_292, n475);
  and g605 (n520, n_292, n518);
  not g606 (n_293, n519);
  not g607 (n_294, n520);
  and g608 (n521, n_293, n_294);
  not g609 (n_295, n521);
  and g610 (n522, n474, n_295);
  not g611 (n_296, n474);
  and g612 (n523, n_296, n_293);
  and g613 (n524, n_294, n523);
  not g614 (n_297, n522);
  not g615 (n_298, n524);
  and g616 (\asquared[13] , n_297, n_298);
  and g617 (n526, \a[9] , \a[13] );
  and g618 (n527, n212, n526);
  and g619 (n528, n209, n484);
  and g620 (n529, \a[3] , \a[13] );
  and g621 (n530, n383, n529);
  not g622 (n_300, n528);
  not g623 (n_301, n530);
  and g624 (n531, n_300, n_301);
  not g625 (n_302, n527);
  not g626 (n_303, n531);
  and g627 (n532, n_302, n_303);
  not g628 (n_304, n532);
  and g629 (n533, \a[3] , n_304);
  and g630 (n534, \a[10] , n533);
  and g631 (n535, n_302, n_304);
  and g632 (n536, \a[0] , \a[13] );
  and g633 (n537, \a[4] , \a[9] );
  not g634 (n_305, n536);
  not g635 (n_306, n537);
  and g636 (n538, n_305, n_306);
  not g637 (n_307, n538);
  and g638 (n539, n535, n_307);
  not g639 (n_308, n534);
  not g640 (n_309, n539);
  and g641 (n540, n_308, n_309);
  not g642 (n_310, n540);
  and g643 (n541, n509, n_310);
  not g644 (n_311, n509);
  and g645 (n542, n_311, n540);
  not g646 (n_312, n541);
  not g647 (n_313, n542);
  and g648 (n543, n_312, n_313);
  and g649 (n544, \a[2] , \a[11] );
  not g650 (n_314, n335);
  not g651 (n_315, n354);
  and g652 (n545, n_314, n_315);
  and g653 (n546, n332, n380);
  not g654 (n_316, n546);
  and g655 (n547, n544, n_316);
  not g656 (n_317, n545);
  and g657 (n548, n_317, n547);
  not g658 (n_318, n548);
  and g659 (n549, n544, n_318);
  and g660 (n550, n_316, n_318);
  and g661 (n551, n_317, n550);
  not g662 (n_319, n549);
  not g663 (n_320, n551);
  and g664 (n552, n_319, n_320);
  not g665 (n_321, n543);
  not g666 (n_322, n552);
  and g667 (n553, n_321, n_322);
  and g668 (n554, n543, n552);
  not g669 (n_323, n553);
  not g670 (n_324, n554);
  and g671 (n555, n_323, n_324);
  and g672 (n556, n_257, n_270);
  not g673 (n_325, \a[12] );
  and g674 (n557, n_325, n503);
  and g675 (n558, \a[12] , n299);
  and g676 (n559, \a[1] , \a[12] );
  not g677 (n_326, \a[7] );
  not g678 (n_327, n559);
  and g679 (n560, n_326, n_327);
  not g680 (n_328, n558);
  not g681 (n_329, n560);
  and g682 (n561, n_328, n_329);
  not g683 (n_330, n561);
  and g684 (n562, n_276, n_330);
  not g685 (n_331, n557);
  not g686 (n_332, n562);
  and g687 (n563, n_331, n_332);
  not g688 (n_333, n489);
  and g689 (n564, n_333, n563);
  not g690 (n_334, n563);
  and g691 (n565, n489, n_334);
  not g692 (n_335, n564);
  not g693 (n_336, n565);
  and g694 (n566, n_335, n_336);
  not g695 (n_337, n566);
  and g696 (n567, n556, n_337);
  not g697 (n_338, n556);
  and g698 (n568, n_338, n566);
  not g699 (n_339, n567);
  not g700 (n_340, n568);
  and g701 (n569, n_339, n_340);
  and g702 (n570, n_285, n_289);
  not g703 (n_341, n569);
  and g704 (n571, n_341, n570);
  not g705 (n_342, n570);
  and g706 (n572, n569, n_342);
  not g707 (n_343, n571);
  not g708 (n_344, n572);
  and g709 (n573, n_343, n_344);
  not g710 (n_345, n555);
  not g711 (n_346, n573);
  and g712 (n574, n_345, n_346);
  and g713 (n575, n555, n573);
  not g714 (n_347, n574);
  not g715 (n_348, n575);
  and g716 (n576, n_347, n_348);
  not g717 (n_349, n523);
  and g718 (n577, n_294, n_349);
  not g719 (n_350, n576);
  and g720 (n578, n_350, n577);
  not g721 (n_351, n577);
  and g722 (n579, n576, n_351);
  not g723 (n_352, n578);
  not g724 (n_353, n579);
  and g725 (\asquared[14] , n_352, n_353);
  and g726 (n581, n_347, n_351);
  not g727 (n_354, n581);
  and g728 (n582, n_348, n_354);
  and g729 (n583, n_340, n_344);
  and g730 (n584, \a[1] , \a[13] );
  not g731 (n_355, n312);
  not g732 (n_356, n584);
  and g733 (n585, n_355, n_356);
  and g734 (n586, n312, n584);
  not g735 (n_357, n550);
  not g736 (n_358, n586);
  and g737 (n587, n_357, n_358);
  not g738 (n_359, n585);
  and g739 (n588, n_359, n587);
  not g740 (n_360, n588);
  and g741 (n589, n_357, n_360);
  and g742 (n590, n_358, n_360);
  and g743 (n591, n_359, n590);
  not g744 (n_361, n589);
  not g745 (n_362, n591);
  and g746 (n592, n_361, n_362);
  not g747 (n_363, n535);
  not g748 (n_364, n592);
  and g749 (n593, n_363, n_364);
  not g750 (n_365, n593);
  and g751 (n594, n_363, n_365);
  and g752 (n595, n_364, n_365);
  not g753 (n_366, n594);
  not g754 (n_367, n595);
  and g755 (n596, n_366, n_367);
  and g756 (n597, n_311, n_310);
  not g757 (n_368, n597);
  and g758 (n598, n_323, n_368);
  and g759 (n599, n596, n598);
  not g760 (n_369, n596);
  not g761 (n_370, n598);
  and g762 (n600, n_369, n_370);
  not g763 (n_371, n599);
  not g764 (n_372, n600);
  and g765 (n601, n_371, n_372);
  and g766 (n602, \a[11] , \a[12] );
  and g767 (n603, n218, n602);
  and g768 (n604, \a[3] , \a[14] );
  and g769 (n605, n449, n604);
  and g770 (n606, \a[12] , \a[14] );
  and g771 (n607, n196, n606);
  not g772 (n_374, n605);
  not g773 (n_375, n607);
  and g774 (n608, n_374, n_375);
  not g775 (n_376, n603);
  not g776 (n_377, n608);
  and g777 (n609, n_376, n_377);
  not g778 (n_378, n609);
  and g779 (n610, n_376, n_378);
  and g780 (n611, \a[2] , \a[12] );
  and g781 (n612, \a[3] , \a[11] );
  not g782 (n_379, n611);
  not g783 (n_380, n612);
  and g784 (n613, n_379, n_380);
  not g785 (n_381, n613);
  and g786 (n614, n610, n_381);
  and g787 (n615, \a[14] , n_378);
  and g788 (n616, \a[0] , n615);
  not g789 (n_382, n614);
  not g790 (n_383, n616);
  and g791 (n617, n_382, n_383);
  and g792 (n618, n226, n484);
  and g793 (n619, \a[4] , \a[10] );
  and g794 (n620, \a[5] , \a[9] );
  not g795 (n_384, n619);
  not g796 (n_385, n620);
  and g797 (n621, n_384, n_385);
  not g798 (n_386, n618);
  not g799 (n_387, n621);
  and g800 (n622, n_386, n_387);
  and g801 (n623, n558, n622);
  not g802 (n_388, n623);
  and g803 (n624, n558, n_388);
  and g804 (n625, n_386, n_388);
  and g805 (n626, n_387, n625);
  not g806 (n_389, n624);
  not g807 (n_390, n626);
  and g808 (n627, n_389, n_390);
  not g809 (n_391, n617);
  not g810 (n_392, n627);
  and g811 (n628, n_391, n_392);
  not g812 (n_393, n628);
  and g813 (n629, n_391, n_393);
  and g814 (n630, n_392, n_393);
  not g815 (n_394, n629);
  not g816 (n_395, n630);
  and g817 (n631, n_394, n_395);
  and g818 (n632, n_331, n_335);
  and g819 (n633, n631, n632);
  not g820 (n_396, n631);
  not g821 (n_397, n632);
  and g822 (n634, n_396, n_397);
  not g823 (n_398, n633);
  not g824 (n_399, n634);
  and g825 (n635, n_398, n_399);
  not g826 (n_400, n635);
  and g827 (n636, n601, n_400);
  not g828 (n_401, n601);
  and g829 (n637, n_401, n635);
  not g830 (n_402, n636);
  not g831 (n_403, n637);
  and g832 (n638, n_402, n_403);
  not g833 (n_404, n583);
  not g834 (n_405, n638);
  and g835 (n639, n_404, n_405);
  and g836 (n640, n583, n638);
  not g837 (n_406, n639);
  not g838 (n_407, n640);
  and g839 (n641, n_406, n_407);
  not g840 (n_408, n641);
  and g841 (n642, n582, n_408);
  not g842 (n_409, n582);
  and g843 (n643, n_409, n_407);
  and g844 (n644, n_406, n643);
  not g845 (n_410, n642);
  not g846 (n_411, n644);
  and g847 (\asquared[15] , n_410, n_411);
  not g848 (n_412, n643);
  and g849 (n646, n_406, n_412);
  and g850 (n647, n601, n635);
  not g851 (n_413, n647);
  and g852 (n648, n_372, n_413);
  and g853 (n649, \a[4] , \a[11] );
  not g854 (n_414, n649);
  and g855 (n650, n_358, n_414);
  and g856 (n651, n586, n649);
  and g857 (n652, \a[1] , \a[14] );
  not g858 (n_415, n652);
  and g859 (n653, \a[8] , n_415);
  not g860 (n_416, \a[8] );
  and g861 (n654, n_416, n652);
  not g862 (n_417, n653);
  not g863 (n_418, n654);
  and g864 (n655, n_417, n_418);
  not g865 (n_419, n651);
  not g866 (n_420, n655);
  and g867 (n656, n_419, n_420);
  not g868 (n_421, n650);
  and g869 (n657, n_421, n656);
  not g870 (n_422, n657);
  and g871 (n658, n_419, n_422);
  and g872 (n659, n_421, n658);
  and g873 (n660, n_420, n_422);
  not g874 (n_423, n659);
  not g875 (n_424, n660);
  and g876 (n661, n_423, n_424);
  and g877 (n662, \a[6] , \a[9] );
  not g878 (n_425, n380);
  not g879 (n_426, n662);
  and g880 (n663, n_425, n_426);
  and g881 (n664, n380, n662);
  not g882 (n_427, n664);
  not g885 (n_428, n663);
  not g887 (n_429, n667);
  and g888 (n668, \a[13] , n_429);
  and g889 (n669, \a[2] , n668);
  and g890 (n670, n_427, n_429);
  and g891 (n671, n_428, n670);
  not g892 (n_430, n669);
  not g893 (n_431, n671);
  and g894 (n672, n_430, n_431);
  not g895 (n_432, n661);
  not g896 (n_433, n672);
  and g897 (n673, n_432, n_433);
  not g898 (n_434, n673);
  and g899 (n674, n_432, n_434);
  and g900 (n675, n_433, n_434);
  not g901 (n_435, n674);
  not g902 (n_436, n675);
  and g903 (n676, n_435, n_436);
  and g904 (n677, n_360, n_365);
  and g905 (n678, n676, n677);
  not g906 (n_437, n676);
  not g907 (n_438, n677);
  and g908 (n679, n_437, n_438);
  not g909 (n_439, n678);
  not g910 (n_440, n679);
  and g911 (n680, n_439, n_440);
  and g912 (n681, n610, n625);
  not g913 (n_441, n610);
  not g914 (n_442, n625);
  and g915 (n682, n_441, n_442);
  not g916 (n_443, n681);
  not g917 (n_444, n682);
  and g918 (n683, n_443, n_444);
  and g919 (n684, \a[5] , \a[10] );
  and g920 (n685, \a[10] , \a[15] );
  and g921 (n686, \a[0] , n685);
  and g922 (n687, \a[3] , n480);
  not g923 (n_446, n686);
  not g924 (n_447, n687);
  and g925 (n688, n_446, n_447);
  and g926 (n689, \a[0] , \a[15] );
  and g927 (n690, \a[3] , \a[12] );
  and g928 (n691, n689, n690);
  not g929 (n_448, n691);
  and g930 (n692, \a[5] , n_448);
  not g931 (n_449, n688);
  and g932 (n693, n_449, n692);
  not g933 (n_450, n693);
  and g934 (n694, n684, n_450);
  and g935 (n695, n_448, n_450);
  not g936 (n_451, n689);
  not g937 (n_452, n690);
  and g938 (n696, n_451, n_452);
  not g939 (n_453, n696);
  and g940 (n697, n695, n_453);
  not g941 (n_454, n694);
  not g942 (n_455, n697);
  and g943 (n698, n_454, n_455);
  not g944 (n_456, n698);
  and g945 (n699, n683, n_456);
  not g946 (n_457, n699);
  and g947 (n700, n683, n_457);
  and g948 (n701, n_456, n_457);
  not g949 (n_458, n700);
  not g950 (n_459, n701);
  and g951 (n702, n_458, n_459);
  and g952 (n703, n_393, n_399);
  and g953 (n704, n702, n703);
  not g954 (n_460, n702);
  not g955 (n_461, n703);
  and g956 (n705, n_460, n_461);
  not g957 (n_462, n704);
  not g958 (n_463, n705);
  and g959 (n706, n_462, n_463);
  not g960 (n_464, n706);
  and g961 (n707, n680, n_464);
  not g962 (n_465, n680);
  and g963 (n708, n_465, n706);
  not g964 (n_466, n707);
  not g965 (n_467, n708);
  and g966 (n709, n_466, n_467);
  not g967 (n_468, n648);
  not g968 (n_469, n709);
  and g969 (n710, n_468, n_469);
  and g970 (n711, n648, n709);
  not g971 (n_470, n710);
  not g972 (n_471, n711);
  and g973 (n712, n_470, n_471);
  not g974 (n_472, n646);
  not g975 (n_473, n712);
  and g976 (n713, n_472, n_473);
  and g977 (n714, n646, n712);
  or g978 (\asquared[16] , n713, n714);
  and g979 (n716, n680, n706);
  not g980 (n_474, n716);
  and g981 (n717, n_463, n_474);
  and g982 (n718, n658, n695);
  not g983 (n_475, n658);
  not g984 (n_476, n695);
  and g985 (n719, n_475, n_476);
  not g986 (n_477, n718);
  not g987 (n_478, n719);
  and g988 (n720, n_477, n_478);
  and g989 (n721, \a[6] , \a[16] );
  and g990 (n722, n383, n721);
  and g991 (n723, \a[10] , \a[11] );
  and g992 (n724, n332, n723);
  and g993 (n725, \a[0] , \a[16] );
  and g994 (n726, n502, n725);
  not g995 (n_480, n724);
  not g996 (n_481, n726);
  and g997 (n727, n_480, n_481);
  not g998 (n_482, n722);
  not g999 (n_483, n727);
  and g1000 (n728, n_482, n_483);
  not g1001 (n_484, n728);
  and g1002 (n729, n502, n_484);
  and g1003 (n730, n_482, n_484);
  and g1004 (n731, \a[6] , \a[10] );
  not g1005 (n_485, n725);
  not g1006 (n_486, n731);
  and g1007 (n732, n_485, n_486);
  not g1008 (n_487, n732);
  and g1009 (n733, n730, n_487);
  not g1010 (n_488, n729);
  not g1011 (n_489, n733);
  and g1012 (n734, n_488, n_489);
  not g1013 (n_490, n734);
  and g1014 (n735, n720, n_490);
  not g1015 (n_491, n735);
  and g1016 (n736, n720, n_491);
  and g1017 (n737, n_490, n_491);
  not g1018 (n_492, n736);
  not g1019 (n_493, n737);
  and g1020 (n738, n_492, n_493);
  and g1021 (n739, n_434, n_440);
  and g1022 (n740, n738, n739);
  not g1023 (n_494, n738);
  not g1024 (n_495, n739);
  and g1025 (n741, n_494, n_495);
  not g1026 (n_496, n740);
  not g1027 (n_497, n741);
  and g1028 (n742, n_496, n_497);
  and g1029 (n743, n_444, n_457);
  and g1030 (n744, \a[4] , \a[12] );
  and g1031 (n745, \a[13] , \a[14] );
  and g1032 (n746, n218, n745);
  and g1033 (n747, n252, n606);
  and g1034 (n748, \a[12] , \a[13] );
  and g1035 (n749, n209, n748);
  not g1036 (n_498, n747);
  not g1037 (n_499, n749);
  and g1038 (n750, n_498, n_499);
  not g1039 (n_500, n746);
  not g1040 (n_501, n750);
  and g1041 (n751, n_500, n_501);
  not g1042 (n_502, n751);
  and g1043 (n752, n744, n_502);
  and g1044 (n753, n_500, n_502);
  and g1045 (n754, \a[2] , \a[14] );
  not g1046 (n_503, n529);
  not g1047 (n_504, n754);
  and g1048 (n755, n_503, n_504);
  not g1049 (n_505, n755);
  and g1050 (n756, n753, n_505);
  not g1051 (n_506, n752);
  not g1052 (n_507, n756);
  and g1053 (n757, n_506, n_507);
  not g1054 (n_508, n743);
  not g1055 (n_509, n757);
  and g1056 (n758, n_508, n_509);
  not g1057 (n_510, n758);
  and g1058 (n759, n_508, n_510);
  and g1059 (n760, n_509, n_510);
  not g1060 (n_511, n759);
  not g1061 (n_512, n760);
  and g1062 (n761, n_511, n_512);
  and g1063 (n762, \a[8] , n652);
  and g1064 (n763, \a[7] , \a[9] );
  and g1065 (n764, \a[1] , \a[15] );
  and g1066 (n765, n763, n764);
  not g1067 (n_513, n763);
  not g1068 (n_514, n764);
  and g1069 (n766, n_513, n_514);
  not g1070 (n_515, n765);
  not g1071 (n_516, n766);
  and g1072 (n767, n_515, n_516);
  and g1073 (n768, n762, n767);
  not g1074 (n_517, n768);
  and g1075 (n769, n762, n_517);
  not g1076 (n_518, n762);
  and g1077 (n770, n_518, n767);
  not g1078 (n_519, n769);
  not g1079 (n_520, n770);
  and g1080 (n771, n_519, n_520);
  not g1081 (n_521, n670);
  not g1082 (n_522, n771);
  and g1083 (n772, n_521, n_522);
  not g1084 (n_523, n772);
  and g1085 (n773, n_521, n_523);
  and g1086 (n774, n_522, n_523);
  not g1087 (n_524, n773);
  not g1088 (n_525, n774);
  and g1089 (n775, n_524, n_525);
  not g1090 (n_526, n761);
  not g1091 (n_527, n775);
  and g1092 (n776, n_526, n_527);
  not g1093 (n_528, n776);
  and g1094 (n777, n_526, n_528);
  and g1095 (n778, n_527, n_528);
  not g1096 (n_529, n777);
  not g1097 (n_530, n778);
  and g1098 (n779, n_529, n_530);
  not g1099 (n_531, n742);
  and g1100 (n780, n_531, n779);
  not g1101 (n_532, n779);
  and g1102 (n781, n742, n_532);
  not g1103 (n_533, n780);
  not g1104 (n_534, n781);
  and g1105 (n782, n_533, n_534);
  not g1106 (n_535, n717);
  and g1107 (n783, n_535, n782);
  not g1108 (n_536, n782);
  and g1109 (n784, n717, n_536);
  not g1110 (n_537, n783);
  not g1111 (n_538, n784);
  and g1112 (n785, n_537, n_538);
  and g1113 (n786, n_472, n_471);
  not g1114 (n_539, n786);
  and g1115 (n787, n_470, n_539);
  not g1116 (n_540, n785);
  and g1117 (n788, n_540, n787);
  not g1118 (n_541, n787);
  and g1119 (n789, n785, n_541);
  not g1120 (n_542, n788);
  not g1121 (n_543, n789);
  and g1122 (\asquared[17] , n_542, n_543);
  and g1123 (n791, n_497, n_534);
  and g1124 (n792, \a[5] , \a[12] );
  and g1125 (n793, \a[0] , \a[17] );
  not g1126 (n_545, n792);
  not g1127 (n_546, n793);
  and g1128 (n794, n_545, n_546);
  and g1129 (n795, n792, n793);
  not g1130 (n_547, n794);
  not g1131 (n_548, n795);
  and g1132 (n796, n_547, n_548);
  and g1133 (n797, n765, n796);
  not g1134 (n_549, n797);
  and g1135 (n798, n_548, n_549);
  and g1136 (n799, n_547, n798);
  and g1137 (n800, n765, n_549);
  not g1138 (n_550, n799);
  not g1139 (n_551, n800);
  and g1140 (n801, n_550, n_551);
  and g1141 (n802, \a[7] , \a[10] );
  not g1142 (n_552, n432);
  not g1143 (n_553, n802);
  and g1144 (n803, n_552, n_553);
  and g1145 (n804, n380, n484);
  not g1146 (n_554, n804);
  and g1147 (n805, n604, n_554);
  not g1148 (n_555, n803);
  and g1149 (n806, n_555, n805);
  not g1150 (n_556, n806);
  and g1151 (n807, n604, n_556);
  and g1152 (n808, n_554, n_556);
  and g1153 (n809, n_555, n808);
  not g1154 (n_557, n807);
  not g1155 (n_558, n809);
  and g1156 (n810, n_557, n_558);
  not g1157 (n_559, n801);
  not g1158 (n_560, n810);
  and g1159 (n811, n_559, n_560);
  not g1160 (n_561, n811);
  and g1161 (n812, n_559, n_561);
  and g1162 (n813, n_560, n_561);
  not g1163 (n_562, n812);
  not g1164 (n_563, n813);
  and g1165 (n814, n_562, n_563);
  and g1166 (n815, \a[6] , \a[11] );
  and g1167 (n816, \a[11] , \a[15] );
  and g1168 (n817, \a[2] , n816);
  and g1169 (n818, \a[11] , \a[13] );
  and g1170 (n819, \a[4] , n818);
  not g1171 (n_564, n817);
  not g1172 (n_565, n819);
  and g1173 (n820, n_564, n_565);
  and g1174 (n821, \a[13] , \a[15] );
  and g1175 (n822, n252, n821);
  not g1176 (n_566, n822);
  and g1177 (n823, \a[6] , n_566);
  not g1178 (n_567, n820);
  and g1179 (n824, n_567, n823);
  not g1180 (n_568, n824);
  and g1181 (n825, n815, n_568);
  and g1182 (n826, n_566, n_568);
  and g1183 (n827, \a[2] , \a[15] );
  and g1184 (n828, \a[4] , \a[13] );
  not g1185 (n_569, n827);
  not g1186 (n_570, n828);
  and g1187 (n829, n_569, n_570);
  not g1188 (n_571, n829);
  and g1189 (n830, n826, n_571);
  not g1190 (n_572, n825);
  not g1191 (n_573, n830);
  and g1192 (n831, n_572, n_573);
  not g1193 (n_574, n814);
  not g1194 (n_575, n831);
  and g1195 (n832, n_574, n_575);
  not g1196 (n_576, n832);
  and g1197 (n833, n_574, n_576);
  and g1198 (n834, n_575, n_576);
  not g1199 (n_577, n833);
  not g1200 (n_578, n834);
  and g1201 (n835, n_577, n_578);
  and g1202 (n836, n_510, n_528);
  and g1203 (n837, n835, n836);
  not g1204 (n_579, n835);
  not g1205 (n_580, n836);
  and g1206 (n838, n_579, n_580);
  not g1207 (n_581, n837);
  not g1208 (n_582, n838);
  and g1209 (n839, n_581, n_582);
  and g1210 (n840, n_517, n_523);
  and g1211 (n841, n_478, n_491);
  and g1212 (n842, n840, n841);
  not g1213 (n_583, n840);
  not g1214 (n_584, n841);
  and g1215 (n843, n_583, n_584);
  not g1216 (n_585, n842);
  not g1217 (n_586, n843);
  and g1218 (n844, n_585, n_586);
  and g1219 (n845, \a[1] , \a[16] );
  not g1220 (n_587, \a[9] );
  not g1221 (n_588, n845);
  and g1222 (n846, n_587, n_588);
  and g1223 (n847, \a[9] , \a[16] );
  and g1224 (n848, \a[1] , n847);
  not g1225 (n_589, n753);
  not g1226 (n_590, n848);
  and g1227 (n849, n_589, n_590);
  not g1228 (n_591, n846);
  and g1229 (n850, n_591, n849);
  not g1230 (n_592, n850);
  and g1231 (n851, n_589, n_592);
  and g1232 (n852, n_590, n_592);
  and g1233 (n853, n_591, n852);
  not g1234 (n_593, n851);
  not g1235 (n_594, n853);
  and g1236 (n854, n_593, n_594);
  not g1237 (n_595, n730);
  not g1238 (n_596, n854);
  and g1239 (n855, n_595, n_596);
  not g1240 (n_597, n855);
  and g1241 (n856, n_595, n_597);
  and g1242 (n857, n_596, n_597);
  not g1243 (n_598, n856);
  not g1244 (n_599, n857);
  and g1245 (n858, n_598, n_599);
  not g1246 (n_600, n844);
  and g1247 (n859, n_600, n858);
  not g1248 (n_601, n858);
  and g1249 (n860, n844, n_601);
  not g1250 (n_602, n859);
  not g1251 (n_603, n860);
  and g1252 (n861, n_602, n_603);
  and g1253 (n862, n839, n861);
  not g1254 (n_604, n839);
  not g1255 (n_605, n861);
  and g1256 (n863, n_604, n_605);
  not g1257 (n_606, n862);
  not g1258 (n_607, n863);
  and g1259 (n864, n_606, n_607);
  not g1260 (n_608, n791);
  and g1261 (n865, n_608, n864);
  not g1262 (n_609, n864);
  and g1263 (n866, n791, n_609);
  not g1264 (n_610, n865);
  not g1265 (n_611, n866);
  and g1266 (n867, n_610, n_611);
  and g1267 (n868, n_538, n_541);
  not g1268 (n_612, n868);
  and g1269 (n869, n_537, n_612);
  not g1270 (n_613, n867);
  and g1271 (n870, n_613, n869);
  not g1272 (n_614, n869);
  and g1273 (n871, n867, n_614);
  not g1274 (n_615, n870);
  not g1275 (n_616, n871);
  and g1276 (\asquared[18] , n_615, n_616);
  and g1277 (n873, n_611, n_614);
  not g1278 (n_617, n873);
  and g1279 (n874, n_610, n_617);
  and g1280 (n875, n_582, n_606);
  and g1281 (n876, \a[7] , \a[18] );
  and g1282 (n877, n449, n876);
  and g1283 (n878, n268, n818);
  not g1284 (n_619, n877);
  not g1285 (n_620, n878);
  and g1286 (n879, n_619, n_620);
  and g1287 (n880, \a[0] , \a[18] );
  and g1288 (n881, \a[5] , \a[13] );
  and g1289 (n882, n880, n881);
  not g1290 (n_621, n879);
  not g1291 (n_622, n882);
  and g1292 (n883, n_621, n_622);
  not g1293 (n_623, n883);
  and g1294 (n884, n_622, n_623);
  not g1295 (n_624, n880);
  not g1296 (n_625, n881);
  and g1297 (n885, n_624, n_625);
  not g1298 (n_626, n885);
  and g1299 (n886, n884, n_626);
  and g1300 (n887, \a[11] , n_623);
  and g1301 (n888, \a[7] , n887);
  not g1302 (n_627, n886);
  not g1303 (n_628, n888);
  and g1304 (n889, n_627, n_628);
  and g1305 (n890, \a[4] , \a[14] );
  and g1306 (n891, \a[15] , \a[16] );
  and g1307 (n892, n218, n891);
  and g1308 (n893, \a[14] , \a[16] );
  and g1309 (n894, n252, n893);
  and g1310 (n895, \a[14] , \a[15] );
  and g1311 (n896, n209, n895);
  not g1312 (n_629, n894);
  not g1313 (n_630, n896);
  and g1314 (n897, n_629, n_630);
  not g1315 (n_631, n892);
  not g1316 (n_632, n897);
  and g1317 (n898, n_631, n_632);
  not g1318 (n_633, n898);
  and g1319 (n899, n890, n_633);
  and g1320 (n900, n_631, n_633);
  and g1321 (n901, \a[3] , \a[15] );
  and g1322 (n902, \a[2] , \a[16] );
  not g1323 (n_634, n901);
  not g1324 (n_635, n902);
  and g1325 (n903, n_634, n_635);
  not g1326 (n_636, n903);
  and g1327 (n904, n900, n_636);
  not g1328 (n_637, n899);
  not g1329 (n_638, n904);
  and g1330 (n905, n_637, n_638);
  not g1331 (n_639, n889);
  not g1332 (n_640, n905);
  and g1333 (n906, n_639, n_640);
  not g1334 (n_641, n906);
  and g1335 (n907, n_639, n_641);
  and g1336 (n908, n_640, n_641);
  not g1337 (n_642, n907);
  not g1338 (n_643, n908);
  and g1339 (n909, n_642, n_643);
  and g1340 (n910, \a[1] , \a[17] );
  and g1341 (n911, n378, n910);
  not g1342 (n_644, n911);
  and g1343 (n912, n378, n_644);
  not g1344 (n_645, n378);
  and g1345 (n913, n_645, n910);
  not g1346 (n_646, n912);
  not g1347 (n_647, n913);
  and g1348 (n914, n_646, n_647);
  and g1349 (n915, \a[6] , \a[12] );
  not g1350 (n_648, n915);
  and g1351 (n916, n_590, n_648);
  and g1352 (n917, n848, n915);
  not g1353 (n_649, n914);
  not g1354 (n_650, n917);
  and g1355 (n918, n_649, n_650);
  not g1356 (n_651, n916);
  and g1357 (n919, n_651, n918);
  not g1358 (n_652, n919);
  and g1359 (n920, n_649, n_652);
  and g1360 (n921, n_650, n_652);
  and g1361 (n922, n_651, n921);
  not g1362 (n_653, n920);
  not g1363 (n_654, n922);
  and g1364 (n923, n_653, n_654);
  not g1365 (n_655, n909);
  not g1366 (n_656, n923);
  and g1367 (n924, n_655, n_656);
  not g1368 (n_657, n924);
  and g1369 (n925, n_655, n_657);
  and g1370 (n926, n_656, n_657);
  not g1371 (n_658, n925);
  not g1372 (n_659, n926);
  and g1373 (n927, n_658, n_659);
  and g1374 (n928, n_586, n_603);
  not g1375 (n_660, n927);
  not g1376 (n_661, n928);
  and g1377 (n929, n_660, n_661);
  not g1378 (n_662, n929);
  and g1379 (n930, n_660, n_662);
  and g1380 (n931, n_661, n_662);
  not g1381 (n_663, n930);
  not g1382 (n_664, n931);
  and g1383 (n932, n_663, n_664);
  and g1384 (n933, n808, n826);
  not g1385 (n_665, n808);
  not g1386 (n_666, n826);
  and g1387 (n934, n_665, n_666);
  not g1388 (n_667, n933);
  not g1389 (n_668, n934);
  and g1390 (n935, n_667, n_668);
  not g1391 (n_669, n935);
  and g1392 (n936, n798, n_669);
  not g1393 (n_670, n798);
  and g1394 (n937, n_670, n935);
  not g1395 (n_671, n936);
  not g1396 (n_672, n937);
  and g1397 (n938, n_671, n_672);
  and g1398 (n939, n_592, n_597);
  and g1399 (n940, n_561, n_576);
  and g1400 (n941, n939, n940);
  not g1401 (n_673, n939);
  not g1402 (n_674, n940);
  and g1403 (n942, n_673, n_674);
  not g1404 (n_675, n941);
  not g1405 (n_676, n942);
  and g1406 (n943, n_675, n_676);
  and g1407 (n944, n938, n943);
  not g1408 (n_677, n938);
  not g1409 (n_678, n943);
  and g1410 (n945, n_677, n_678);
  not g1411 (n_679, n944);
  not g1412 (n_680, n945);
  and g1413 (n946, n_679, n_680);
  not g1414 (n_681, n932);
  and g1415 (n947, n_681, n946);
  not g1416 (n_682, n946);
  and g1417 (n948, n932, n_682);
  not g1418 (n_683, n947);
  not g1419 (n_684, n948);
  and g1420 (n949, n_683, n_684);
  not g1421 (n_685, n875);
  and g1422 (n950, n_685, n949);
  not g1423 (n_686, n949);
  and g1424 (n951, n875, n_686);
  not g1425 (n_687, n950);
  not g1426 (n_688, n951);
  and g1427 (n952, n_687, n_688);
  not g1428 (n_689, n952);
  and g1429 (n953, n874, n_689);
  not g1430 (n_690, n874);
  and g1431 (n954, n_690, n_688);
  and g1432 (n955, n_687, n954);
  not g1433 (n_691, n953);
  not g1434 (n_692, n955);
  and g1435 (\asquared[19] , n_691, n_692);
  and g1436 (n957, n884, n921);
  not g1437 (n_693, n884);
  not g1438 (n_694, n921);
  and g1439 (n958, n_693, n_694);
  not g1440 (n_695, n957);
  not g1441 (n_696, n958);
  and g1442 (n959, n_695, n_696);
  and g1443 (n960, \a[3] , \a[16] );
  and g1444 (n961, \a[8] , \a[11] );
  not g1445 (n_697, n484);
  not g1446 (n_698, n961);
  and g1447 (n962, n_697, n_698);
  and g1448 (n963, n484, n961);
  not g1449 (n_699, n963);
  and g1450 (n964, n960, n_699);
  not g1451 (n_700, n962);
  and g1452 (n965, n_700, n964);
  not g1453 (n_701, n965);
  and g1454 (n966, n960, n_701);
  and g1455 (n967, n_699, n_701);
  and g1456 (n968, n_700, n967);
  not g1457 (n_702, n966);
  not g1458 (n_703, n968);
  and g1459 (n969, n_702, n_703);
  not g1460 (n_704, n969);
  and g1461 (n970, n959, n_704);
  not g1462 (n_705, n970);
  and g1463 (n971, n959, n_705);
  and g1464 (n972, n_704, n_705);
  not g1465 (n_706, n971);
  not g1466 (n_707, n972);
  and g1467 (n973, n_706, n_707);
  and g1468 (n974, n_641, n_657);
  and g1469 (n975, \a[1] , \a[18] );
  not g1470 (n_708, n975);
  and g1471 (n976, n911, n_708);
  not g1472 (n_709, n976);
  and g1473 (n977, n911, n_709);
  not g1474 (n_710, \a[10] );
  and g1475 (n978, n_710, n_708);
  and g1476 (n979, \a[10] , n975);
  not g1477 (n_711, n979);
  and g1478 (n980, n_709, n_711);
  not g1479 (n_712, n978);
  and g1480 (n981, n_712, n980);
  not g1481 (n_713, n977);
  not g1482 (n_714, n981);
  and g1483 (n982, n_713, n_714);
  not g1484 (n_715, n900);
  not g1485 (n_716, n982);
  and g1486 (n983, n_715, n_716);
  and g1487 (n984, n900, n_714);
  and g1488 (n985, n_713, n984);
  not g1489 (n_717, n983);
  not g1490 (n_718, n985);
  and g1491 (n986, n_717, n_718);
  not g1492 (n_719, n974);
  and g1493 (n987, n_719, n986);
  not g1494 (n_720, n986);
  and g1495 (n988, n974, n_720);
  not g1496 (n_721, n987);
  not g1497 (n_722, n988);
  and g1498 (n989, n_721, n_722);
  not g1499 (n_723, n973);
  and g1500 (n990, n_723, n989);
  not g1501 (n_724, n989);
  and g1502 (n991, n973, n_724);
  not g1503 (n_725, n990);
  not g1504 (n_726, n991);
  and g1505 (n992, n_725, n_726);
  and g1506 (n993, \a[15] , \a[17] );
  and g1507 (n994, n252, n993);
  and g1508 (n995, \a[15] , n212);
  and g1509 (n996, \a[17] , n196);
  not g1510 (n_727, n995);
  not g1511 (n_728, n996);
  and g1512 (n997, n_727, n_728);
  not g1513 (n_730, n994);
  and g1514 (n998, \a[19] , n_730);
  not g1515 (n_731, n997);
  and g1516 (n999, n_731, n998);
  not g1517 (n_732, n999);
  and g1518 (n1000, n_730, n_732);
  and g1519 (n1001, \a[2] , \a[17] );
  and g1520 (n1002, \a[4] , \a[15] );
  not g1521 (n_733, n1001);
  not g1522 (n_734, n1002);
  and g1523 (n1003, n_733, n_734);
  not g1524 (n_735, n1003);
  and g1525 (n1004, n1000, n_735);
  and g1526 (n1005, \a[19] , n_732);
  and g1527 (n1006, \a[0] , n1005);
  not g1528 (n_736, n1004);
  not g1529 (n_737, n1006);
  and g1530 (n1007, n_736, n_737);
  and g1531 (n1008, n335, n748);
  and g1532 (n1009, n268, n606);
  and g1533 (n1010, n332, n745);
  not g1534 (n_738, n1009);
  not g1535 (n_739, n1010);
  and g1536 (n1011, n_738, n_739);
  not g1537 (n_740, n1008);
  not g1538 (n_741, n1011);
  and g1539 (n1012, n_740, n_741);
  not g1540 (n_742, n1012);
  and g1541 (n1013, \a[14] , n_742);
  and g1542 (n1014, \a[5] , n1013);
  and g1543 (n1015, n_740, n_742);
  and g1544 (n1016, \a[6] , \a[13] );
  and g1545 (n1017, \a[7] , \a[12] );
  not g1546 (n_743, n1016);
  not g1547 (n_744, n1017);
  and g1548 (n1018, n_743, n_744);
  not g1549 (n_745, n1018);
  and g1550 (n1019, n1015, n_745);
  not g1551 (n_746, n1014);
  not g1552 (n_747, n1019);
  and g1553 (n1020, n_746, n_747);
  not g1554 (n_748, n1007);
  not g1555 (n_749, n1020);
  and g1556 (n1021, n_748, n_749);
  not g1557 (n_750, n1021);
  and g1558 (n1022, n_748, n_750);
  and g1559 (n1023, n_749, n_750);
  not g1560 (n_751, n1022);
  not g1561 (n_752, n1023);
  and g1562 (n1024, n_751, n_752);
  and g1563 (n1025, n_668, n_672);
  and g1564 (n1026, n1024, n1025);
  not g1565 (n_753, n1024);
  not g1566 (n_754, n1025);
  and g1567 (n1027, n_753, n_754);
  not g1568 (n_755, n1026);
  not g1569 (n_756, n1027);
  and g1570 (n1028, n_755, n_756);
  and g1571 (n1029, n_676, n_679);
  not g1572 (n_757, n1029);
  and g1573 (n1030, n1028, n_757);
  not g1574 (n_758, n1028);
  and g1575 (n1031, n_758, n1029);
  not g1576 (n_759, n1030);
  not g1577 (n_760, n1031);
  and g1578 (n1032, n_759, n_760);
  and g1579 (n1033, n992, n1032);
  not g1580 (n_761, n992);
  not g1581 (n_762, n1032);
  and g1582 (n1034, n_761, n_762);
  not g1583 (n_763, n1033);
  not g1584 (n_764, n1034);
  and g1585 (n1035, n_763, n_764);
  and g1586 (n1036, n_662, n_683);
  not g1587 (n_765, n1035);
  and g1588 (n1037, n_765, n1036);
  not g1589 (n_766, n1036);
  and g1590 (n1038, n1035, n_766);
  not g1591 (n_767, n1037);
  not g1592 (n_768, n1038);
  and g1593 (n1039, n_767, n_768);
  not g1594 (n_769, n954);
  and g1595 (n1040, n_687, n_769);
  not g1596 (n_770, n1039);
  and g1597 (n1041, n_770, n1040);
  not g1598 (n_771, n1040);
  and g1599 (n1042, n1039, n_771);
  not g1600 (n_772, n1041);
  not g1601 (n_773, n1042);
  and g1602 (\asquared[20] , n_772, n_773);
  and g1603 (n1044, n_767, n_771);
  not g1604 (n_774, n1044);
  and g1605 (n1045, n_768, n_774);
  and g1606 (n1046, n_759, n_763);
  and g1607 (n1047, n_709, n_717);
  and g1608 (n1048, \a[16] , \a[17] );
  and g1609 (n1049, n209, n1048);
  and g1610 (n1050, \a[16] , \a[18] );
  and g1611 (n1051, n252, n1050);
  and g1612 (n1052, \a[17] , \a[18] );
  and g1613 (n1053, n218, n1052);
  not g1614 (n_775, n1051);
  not g1615 (n_776, n1053);
  and g1616 (n1054, n_775, n_776);
  not g1617 (n_777, n1049);
  not g1618 (n_778, n1054);
  and g1619 (n1055, n_777, n_778);
  not g1620 (n_779, n1055);
  and g1621 (n1056, \a[18] , n_779);
  and g1622 (n1057, \a[2] , n1056);
  and g1623 (n1058, n_777, n_779);
  and g1624 (n1059, \a[3] , \a[17] );
  and g1625 (n1060, \a[4] , \a[16] );
  not g1626 (n_780, n1059);
  not g1627 (n_781, n1060);
  and g1628 (n1061, n_780, n_781);
  not g1629 (n_782, n1061);
  and g1630 (n1062, n1058, n_782);
  not g1631 (n_783, n1057);
  not g1632 (n_784, n1062);
  and g1633 (n1063, n_783, n_784);
  not g1634 (n_785, n1047);
  not g1635 (n_786, n1063);
  and g1636 (n1064, n_785, n_786);
  not g1637 (n_787, n1064);
  and g1638 (n1065, n_785, n_787);
  and g1639 (n1066, n_786, n_787);
  not g1640 (n_788, n1065);
  not g1641 (n_789, n1066);
  and g1642 (n1067, n_788, n_789);
  and g1643 (n1068, n_696, n_705);
  and g1644 (n1069, n1067, n1068);
  not g1645 (n_790, n1067);
  not g1646 (n_791, n1068);
  and g1647 (n1070, n_790, n_791);
  not g1648 (n_792, n1069);
  not g1649 (n_793, n1070);
  and g1650 (n1071, n_792, n_793);
  and g1651 (n1072, n_721, n_725);
  not g1652 (n_794, n1071);
  and g1653 (n1073, n_794, n1072);
  not g1654 (n_795, n1072);
  and g1655 (n1074, n1071, n_795);
  not g1656 (n_796, n1073);
  not g1657 (n_797, n1074);
  and g1658 (n1075, n_796, n_797);
  and g1659 (n1076, \a[9] , \a[11] );
  and g1660 (n1077, \a[1] , \a[19] );
  not g1661 (n_798, n1076);
  not g1662 (n_799, n1077);
  and g1663 (n1078, n_798, n_799);
  and g1664 (n1079, n1076, n1077);
  not g1665 (n_800, n967);
  not g1666 (n_801, n1079);
  and g1667 (n1080, n_800, n_801);
  not g1668 (n_802, n1078);
  and g1669 (n1081, n_802, n1080);
  not g1670 (n_803, n1081);
  and g1671 (n1082, n_800, n_803);
  and g1672 (n1083, n_801, n_803);
  and g1673 (n1084, n_802, n1083);
  not g1674 (n_804, n1082);
  not g1675 (n_805, n1084);
  and g1676 (n1085, n_804, n_805);
  not g1677 (n_806, n1000);
  not g1678 (n_807, n1085);
  and g1679 (n1086, n_806, n_807);
  not g1680 (n_808, n1086);
  and g1681 (n1087, n_806, n_808);
  and g1682 (n1088, n_807, n_808);
  not g1683 (n_809, n1087);
  not g1684 (n_810, n1088);
  and g1685 (n1089, n_809, n_810);
  and g1686 (n1090, n_750, n_756);
  and g1687 (n1091, n1089, n1090);
  not g1688 (n_811, n1089);
  not g1689 (n_812, n1090);
  and g1690 (n1092, n_811, n_812);
  not g1691 (n_813, n1091);
  not g1692 (n_814, n1092);
  and g1693 (n1093, n_813, n_814);
  and g1694 (n1094, \a[0] , \a[20] );
  and g1695 (n1095, \a[7] , \a[13] );
  not g1696 (n_816, n1094);
  not g1697 (n_817, n1095);
  and g1698 (n1096, n_816, n_817);
  and g1699 (n1097, n1094, n1095);
  not g1700 (n_818, n1096);
  not g1701 (n_819, n1097);
  and g1702 (n1098, n_818, n_819);
  and g1703 (n1099, n979, n1098);
  not g1704 (n_820, n1098);
  and g1705 (n1100, n_711, n_820);
  not g1706 (n_821, n1099);
  not g1707 (n_822, n1100);
  and g1708 (n1101, n_821, n_822);
  not g1709 (n_823, n1015);
  and g1710 (n1102, n_823, n1101);
  not g1711 (n_824, n1101);
  and g1712 (n1103, n1015, n_824);
  not g1713 (n_825, n1102);
  not g1714 (n_826, n1103);
  and g1715 (n1104, n_825, n_826);
  and g1716 (n1105, n332, n895);
  and g1717 (n1106, n312, n606);
  and g1718 (n1107, \a[8] , \a[15] );
  and g1719 (n1108, n792, n1107);
  not g1720 (n_827, n1106);
  not g1721 (n_828, n1108);
  and g1722 (n1109, n_827, n_828);
  not g1723 (n_829, n1105);
  not g1724 (n_830, n1109);
  and g1725 (n1110, n_829, n_830);
  not g1726 (n_831, n1110);
  and g1727 (n1111, \a[12] , n_831);
  and g1728 (n1112, \a[8] , n1111);
  and g1729 (n1113, n_829, n_831);
  and g1730 (n1114, \a[5] , \a[15] );
  and g1731 (n1115, \a[6] , \a[14] );
  not g1732 (n_832, n1114);
  not g1733 (n_833, n1115);
  and g1734 (n1116, n_832, n_833);
  not g1735 (n_834, n1116);
  and g1736 (n1117, n1113, n_834);
  not g1737 (n_835, n1112);
  not g1738 (n_836, n1117);
  and g1739 (n1118, n_835, n_836);
  not g1740 (n_837, n1118);
  and g1741 (n1119, n1104, n_837);
  not g1742 (n_838, n1119);
  and g1743 (n1120, n1104, n_838);
  and g1744 (n1121, n_837, n_838);
  not g1745 (n_839, n1120);
  not g1746 (n_840, n1121);
  and g1747 (n1122, n_839, n_840);
  not g1748 (n_841, n1122);
  and g1749 (n1123, n1093, n_841);
  not g1750 (n_842, n1093);
  and g1751 (n1124, n_842, n1122);
  not g1752 (n_843, n1124);
  and g1753 (n1125, n1075, n_843);
  not g1754 (n_844, n1123);
  and g1755 (n1126, n_844, n1125);
  not g1756 (n_845, n1126);
  and g1757 (n1127, n1075, n_845);
  and g1758 (n1128, n_843, n_845);
  and g1759 (n1129, n_844, n1128);
  not g1760 (n_846, n1127);
  not g1761 (n_847, n1129);
  and g1762 (n1130, n_846, n_847);
  not g1763 (n_848, n1046);
  not g1764 (n_849, n1130);
  and g1765 (n1131, n_848, n_849);
  and g1766 (n1132, n1046, n1130);
  not g1767 (n_850, n1131);
  not g1768 (n_851, n1132);
  and g1769 (n1133, n_850, n_851);
  not g1770 (n_852, n1045);
  and g1771 (n1134, n_852, n1133);
  not g1772 (n_853, n1133);
  and g1773 (n1135, n1045, n_853);
  not g1774 (n_854, n1134);
  not g1775 (n_855, n1135);
  and g1776 (\asquared[21] , n_854, n_855);
  and g1777 (n1137, n_797, n_845);
  and g1778 (n1138, n1058, n1113);
  not g1779 (n_856, n1058);
  not g1780 (n_857, n1113);
  and g1781 (n1139, n_856, n_857);
  not g1782 (n_858, n1138);
  not g1783 (n_859, n1139);
  and g1784 (n1140, n_858, n_859);
  and g1785 (n1141, n_819, n_821);
  not g1786 (n_860, n1140);
  and g1787 (n1142, n_860, n1141);
  not g1788 (n_861, n1141);
  and g1789 (n1143, n1140, n_861);
  not g1790 (n_862, n1142);
  not g1791 (n_863, n1143);
  and g1792 (n1144, n_862, n_863);
  and g1793 (n1145, n_787, n_793);
  not g1794 (n_864, n1144);
  and g1795 (n1146, n_864, n1145);
  not g1796 (n_865, n1145);
  and g1797 (n1147, n1144, n_865);
  not g1798 (n_866, n1146);
  not g1799 (n_867, n1147);
  and g1800 (n1148, n_866, n_867);
  and g1801 (n1149, \a[18] , \a[19] );
  and g1802 (n1150, n218, n1149);
  and g1803 (n1151, \a[19] , n902);
  and g1804 (n1152, \a[3] , n1050);
  not g1805 (n_868, n1151);
  not g1806 (n_869, n1152);
  and g1807 (n1153, n_868, n_869);
  not g1808 (n_870, n1150);
  and g1809 (n1154, \a[5] , n_870);
  not g1810 (n_871, n1153);
  and g1811 (n1155, n_871, n1154);
  not g1812 (n_872, n1155);
  and g1813 (n1156, n_870, n_872);
  and g1814 (n1157, \a[2] , \a[19] );
  and g1815 (n1158, \a[3] , \a[18] );
  not g1816 (n_873, n1157);
  not g1817 (n_874, n1158);
  and g1818 (n1159, n_873, n_874);
  not g1819 (n_875, n1159);
  and g1820 (n1160, n1156, n_875);
  and g1821 (n1161, \a[16] , n_872);
  and g1822 (n1162, \a[5] , n1161);
  not g1823 (n_876, n1160);
  not g1824 (n_877, n1162);
  and g1825 (n1163, n_876, n_877);
  and g1826 (n1164, n380, n745);
  and g1827 (n1165, n312, n821);
  and g1828 (n1166, n335, n895);
  not g1829 (n_878, n1165);
  not g1830 (n_879, n1166);
  and g1831 (n1167, n_878, n_879);
  not g1832 (n_880, n1164);
  not g1833 (n_881, n1167);
  and g1834 (n1168, n_880, n_881);
  not g1835 (n_882, n1168);
  and g1836 (n1169, \a[15] , n_882);
  and g1837 (n1170, \a[6] , n1169);
  and g1838 (n1171, n_880, n_882);
  and g1839 (n1172, \a[7] , \a[14] );
  and g1840 (n1173, \a[8] , \a[13] );
  not g1841 (n_883, n1172);
  not g1842 (n_884, n1173);
  and g1843 (n1174, n_883, n_884);
  not g1844 (n_885, n1174);
  and g1845 (n1175, n1171, n_885);
  not g1846 (n_886, n1170);
  not g1847 (n_887, n1175);
  and g1848 (n1176, n_886, n_887);
  not g1849 (n_888, n1163);
  not g1850 (n_889, n1176);
  and g1851 (n1177, n_888, n_889);
  not g1852 (n_890, n1177);
  and g1853 (n1178, n_888, n_890);
  and g1854 (n1179, n_889, n_890);
  not g1855 (n_891, n1178);
  not g1856 (n_892, n1179);
  and g1857 (n1180, n_891, n_892);
  and g1858 (n1181, \a[4] , \a[17] );
  and g1859 (n1182, \a[9] , \a[12] );
  not g1860 (n_893, n723);
  not g1861 (n_894, n1182);
  and g1862 (n1183, n_893, n_894);
  and g1863 (n1184, n484, n602);
  not g1864 (n_895, n1184);
  and g1865 (n1185, n1181, n_895);
  not g1866 (n_896, n1183);
  and g1867 (n1186, n_896, n1185);
  not g1868 (n_897, n1186);
  and g1869 (n1187, n1181, n_897);
  and g1870 (n1188, n_895, n_897);
  and g1871 (n1189, n_896, n1188);
  not g1872 (n_898, n1187);
  not g1873 (n_899, n1189);
  and g1874 (n1190, n_898, n_899);
  not g1875 (n_900, n1180);
  not g1876 (n_901, n1190);
  and g1877 (n1191, n_900, n_901);
  not g1878 (n_902, n1191);
  and g1879 (n1192, n_900, n_902);
  and g1880 (n1193, n_901, n_902);
  not g1881 (n_903, n1192);
  not g1882 (n_904, n1193);
  and g1883 (n1194, n_903, n_904);
  not g1884 (n_905, n1148);
  and g1885 (n1195, n_905, n1194);
  not g1886 (n_906, n1194);
  and g1887 (n1196, n1148, n_906);
  not g1888 (n_907, n1195);
  not g1889 (n_908, n1196);
  and g1890 (n1197, n_907, n_908);
  and g1891 (n1198, n_803, n_808);
  and g1892 (n1199, \a[0] , \a[21] );
  not g1893 (n_910, n1199);
  and g1894 (n1200, n1079, n_910);
  and g1895 (n1201, n_801, n1199);
  not g1896 (n_911, n1200);
  not g1897 (n_912, n1201);
  and g1898 (n1202, n_911, n_912);
  and g1899 (n1203, \a[1] , \a[20] );
  and g1900 (n1204, \a[11] , n1203);
  not g1901 (n_913, n1204);
  and g1902 (n1205, \a[11] , n_913);
  and g1903 (n1206, n1203, n_913);
  not g1904 (n_914, n1205);
  not g1905 (n_915, n1206);
  and g1906 (n1207, n_914, n_915);
  not g1907 (n_916, n1202);
  not g1908 (n_917, n1207);
  and g1909 (n1208, n_916, n_917);
  and g1910 (n1209, n1202, n1207);
  not g1911 (n_918, n1208);
  not g1912 (n_919, n1209);
  and g1913 (n1210, n_918, n_919);
  not g1914 (n_920, n1210);
  and g1915 (n1211, n1198, n_920);
  not g1916 (n_921, n1198);
  and g1917 (n1212, n_921, n1210);
  not g1918 (n_922, n1211);
  not g1919 (n_923, n1212);
  and g1920 (n1213, n_922, n_923);
  and g1921 (n1214, n_825, n_838);
  not g1922 (n_924, n1213);
  and g1923 (n1215, n_924, n1214);
  not g1924 (n_925, n1214);
  and g1925 (n1216, n1213, n_925);
  not g1926 (n_926, n1215);
  not g1927 (n_927, n1216);
  and g1928 (n1217, n_926, n_927);
  and g1929 (n1218, n_814, n_844);
  not g1930 (n_928, n1218);
  and g1931 (n1219, n1217, n_928);
  not g1932 (n_929, n1217);
  and g1933 (n1220, n_929, n1218);
  not g1934 (n_930, n1219);
  not g1935 (n_931, n1220);
  and g1936 (n1221, n_930, n_931);
  and g1937 (n1222, n1197, n1221);
  not g1938 (n_932, n1197);
  not g1939 (n_933, n1221);
  and g1940 (n1223, n_932, n_933);
  not g1941 (n_934, n1222);
  not g1942 (n_935, n1223);
  and g1943 (n1224, n_934, n_935);
  not g1944 (n_936, n1137);
  and g1945 (n1225, n_936, n1224);
  not g1946 (n_937, n1224);
  and g1947 (n1226, n1137, n_937);
  not g1948 (n_938, n1225);
  not g1949 (n_939, n1226);
  and g1950 (n1227, n_938, n_939);
  and g1951 (n1228, n_852, n_851);
  not g1952 (n_940, n1228);
  and g1953 (n1229, n_850, n_940);
  not g1954 (n_941, n1227);
  and g1955 (n1230, n_941, n1229);
  not g1956 (n_942, n1229);
  and g1957 (n1231, n1227, n_942);
  not g1958 (n_943, n1230);
  not g1959 (n_944, n1231);
  and g1960 (\asquared[22] , n_943, n_944);
  and g1961 (n1233, n_939, n_942);
  not g1962 (n_945, n1233);
  and g1963 (n1234, n_938, n_945);
  and g1964 (n1235, n_930, n_934);
  and g1965 (n1236, n1156, n1171);
  not g1966 (n_946, n1156);
  not g1967 (n_947, n1171);
  and g1968 (n1237, n_946, n_947);
  not g1969 (n_948, n1236);
  not g1970 (n_949, n1237);
  and g1971 (n1238, n_948, n_949);
  and g1972 (n1239, n1079, n1199);
  not g1973 (n_950, n1239);
  and g1974 (n1240, n_918, n_950);
  not g1975 (n_951, n1238);
  and g1976 (n1241, n_951, n1240);
  not g1977 (n_952, n1240);
  and g1978 (n1242, n1238, n_952);
  not g1979 (n_953, n1241);
  not g1980 (n_954, n1242);
  and g1981 (n1243, n_953, n_954);
  and g1982 (n1244, n_923, n_927);
  not g1983 (n_955, n1243);
  and g1984 (n1245, n_955, n1244);
  not g1985 (n_956, n1244);
  and g1986 (n1246, n1243, n_956);
  not g1987 (n_957, n1245);
  not g1988 (n_958, n1246);
  and g1989 (n1247, n_957, n_958);
  and g1990 (n1248, \a[7] , \a[15] );
  and g1991 (n1249, \a[8] , \a[14] );
  not g1992 (n_959, n1248);
  not g1993 (n_960, n1249);
  and g1994 (n1250, n_959, n_960);
  and g1995 (n1251, n380, n895);
  not g1996 (n_961, n1251);
  not g1999 (n_963, n1250);
  not g2001 (n_964, n1254);
  and g2002 (n1255, n_961, n_964);
  and g2003 (n1256, n_963, n1255);
  and g2004 (n1257, \a[22] , n_964);
  and g2005 (n1258, \a[0] , n1257);
  not g2006 (n_965, n1256);
  not g2007 (n_966, n1258);
  and g2008 (n1259, n_965, n_966);
  and g2009 (n1260, \a[2] , \a[20] );
  not g2010 (n_967, n721);
  not g2011 (n_968, n1260);
  and g2012 (n1261, n_967, n_968);
  and g2013 (n1262, n721, n1260);
  not g2014 (n_969, n1262);
  and g2015 (n1263, n526, n_969);
  not g2016 (n_970, n1261);
  and g2017 (n1264, n_970, n1263);
  not g2018 (n_971, n1264);
  and g2019 (n1265, n526, n_971);
  and g2020 (n1266, n_969, n_971);
  and g2021 (n1267, n_970, n1266);
  not g2022 (n_972, n1265);
  not g2023 (n_973, n1267);
  and g2024 (n1268, n_972, n_973);
  not g2025 (n_974, n1259);
  not g2026 (n_975, n1268);
  and g2027 (n1269, n_974, n_975);
  not g2028 (n_976, n1269);
  and g2029 (n1270, n_974, n_976);
  and g2030 (n1271, n_975, n_976);
  not g2031 (n_977, n1270);
  not g2032 (n_978, n1271);
  and g2033 (n1272, n_977, n_978);
  and g2034 (n1273, \a[3] , \a[19] );
  and g2035 (n1274, n226, n1052);
  and g2036 (n1275, n209, n1149);
  and g2037 (n1276, \a[5] , \a[17] );
  and g2038 (n1277, n1273, n1276);
  not g2039 (n_979, n1275);
  not g2040 (n_980, n1277);
  and g2041 (n1278, n_979, n_980);
  not g2042 (n_981, n1274);
  not g2043 (n_982, n1278);
  and g2044 (n1279, n_981, n_982);
  not g2045 (n_983, n1279);
  and g2046 (n1280, n1273, n_983);
  and g2047 (n1281, n_981, n_983);
  and g2048 (n1282, \a[4] , \a[18] );
  not g2049 (n_984, n1276);
  not g2050 (n_985, n1282);
  and g2051 (n1283, n_984, n_985);
  not g2052 (n_986, n1283);
  and g2053 (n1284, n1281, n_986);
  not g2054 (n_987, n1280);
  not g2055 (n_988, n1284);
  and g2056 (n1285, n_987, n_988);
  not g2057 (n_989, n1272);
  not g2058 (n_990, n1285);
  and g2059 (n1286, n_989, n_990);
  not g2060 (n_991, n1286);
  and g2061 (n1287, n_989, n_991);
  and g2062 (n1288, n_990, n_991);
  not g2063 (n_992, n1287);
  not g2064 (n_993, n1288);
  and g2065 (n1289, n_992, n_993);
  not g2066 (n_994, n1247);
  and g2067 (n1290, n_994, n1289);
  not g2068 (n_995, n1289);
  and g2069 (n1291, n1247, n_995);
  not g2070 (n_996, n1290);
  not g2071 (n_997, n1291);
  and g2072 (n1292, n_996, n_997);
  and g2073 (n1293, n_867, n_908);
  and g2074 (n1294, n_890, n_902);
  and g2075 (n1295, n_859, n_863);
  and g2076 (n1296, \a[1] , \a[21] );
  and g2077 (n1297, n480, n1296);
  not g2078 (n_998, n480);
  not g2079 (n_999, n1296);
  and g2080 (n1298, n_998, n_999);
  not g2081 (n_1000, n1297);
  not g2082 (n_1001, n1298);
  and g2083 (n1299, n_1000, n_1001);
  and g2084 (n1300, n1204, n1299);
  not g2085 (n_1002, n1299);
  and g2086 (n1301, n_913, n_1002);
  not g2087 (n_1003, n1300);
  not g2088 (n_1004, n1301);
  and g2089 (n1302, n_1003, n_1004);
  not g2090 (n_1005, n1188);
  and g2091 (n1303, n_1005, n1302);
  not g2092 (n_1006, n1302);
  and g2093 (n1304, n1188, n_1006);
  not g2094 (n_1007, n1303);
  not g2095 (n_1008, n1304);
  and g2096 (n1305, n_1007, n_1008);
  not g2097 (n_1009, n1295);
  and g2098 (n1306, n_1009, n1305);
  not g2099 (n_1010, n1306);
  and g2100 (n1307, n_1009, n_1010);
  and g2101 (n1308, n1305, n_1010);
  not g2102 (n_1011, n1307);
  not g2103 (n_1012, n1308);
  and g2104 (n1309, n_1011, n_1012);
  not g2105 (n_1013, n1294);
  not g2106 (n_1014, n1309);
  and g2107 (n1310, n_1013, n_1014);
  and g2108 (n1311, n1294, n_1012);
  and g2109 (n1312, n_1011, n1311);
  not g2110 (n_1015, n1310);
  not g2111 (n_1016, n1312);
  and g2112 (n1313, n_1015, n_1016);
  not g2113 (n_1017, n1293);
  and g2114 (n1314, n_1017, n1313);
  not g2115 (n_1018, n1314);
  and g2116 (n1315, n_1017, n_1018);
  and g2117 (n1316, n1313, n_1018);
  not g2118 (n_1019, n1315);
  not g2119 (n_1020, n1316);
  and g2120 (n1317, n_1019, n_1020);
  not g2121 (n_1021, n1317);
  and g2122 (n1318, n1292, n_1021);
  not g2123 (n_1022, n1292);
  and g2124 (n1319, n_1022, n_1020);
  and g2125 (n1320, n_1019, n1319);
  not g2126 (n_1023, n1318);
  not g2127 (n_1024, n1320);
  and g2128 (n1321, n_1023, n_1024);
  not g2129 (n_1025, n1235);
  and g2130 (n1322, n_1025, n1321);
  not g2131 (n_1026, n1321);
  and g2132 (n1323, n1235, n_1026);
  not g2133 (n_1027, n1322);
  not g2134 (n_1028, n1323);
  and g2135 (n1324, n_1027, n_1028);
  not g2136 (n_1029, n1324);
  and g2137 (n1325, n1234, n_1029);
  not g2138 (n_1030, n1234);
  and g2139 (n1326, n_1030, n_1028);
  and g2140 (n1327, n_1027, n1326);
  not g2141 (n_1031, n1325);
  not g2142 (n_1032, n1327);
  and g2143 (\asquared[23] , n_1031, n_1032);
  and g2144 (n1329, n_1018, n_1023);
  and g2145 (n1330, n_1010, n_1015);
  and g2146 (n1331, \a[18] , \a[20] );
  and g2147 (n1332, n300, n1331);
  and g2148 (n1333, \a[17] , \a[20] );
  and g2149 (n1334, n340, n1333);
  and g2150 (n1335, n332, n1052);
  not g2151 (n_1033, n1334);
  not g2152 (n_1034, n1335);
  and g2153 (n1336, n_1033, n_1034);
  not g2154 (n_1035, n1332);
  not g2155 (n_1036, n1336);
  and g2156 (n1337, n_1035, n_1036);
  not g2157 (n_1037, n1337);
  and g2158 (n1338, n_1035, n_1037);
  and g2159 (n1339, \a[3] , \a[20] );
  and g2160 (n1340, \a[5] , \a[18] );
  not g2161 (n_1038, n1339);
  not g2162 (n_1039, n1340);
  and g2163 (n1341, n_1038, n_1039);
  not g2164 (n_1040, n1341);
  and g2165 (n1342, n1338, n_1040);
  and g2166 (n1343, \a[17] , n_1037);
  and g2167 (n1344, \a[6] , n1343);
  not g2168 (n_1041, n1342);
  not g2169 (n_1042, n1344);
  and g2170 (n1345, n_1041, n_1042);
  and g2171 (n1346, \a[4] , \a[19] );
  and g2172 (n1347, \a[10] , \a[13] );
  not g2173 (n_1043, n602);
  not g2174 (n_1044, n1347);
  and g2175 (n1348, n_1043, n_1044);
  and g2176 (n1349, n723, n748);
  not g2177 (n_1045, n1349);
  and g2178 (n1350, n1346, n_1045);
  not g2179 (n_1046, n1348);
  and g2180 (n1351, n_1046, n1350);
  not g2181 (n_1047, n1351);
  and g2182 (n1352, n1346, n_1047);
  and g2183 (n1353, n_1045, n_1047);
  and g2184 (n1354, n_1046, n1353);
  not g2185 (n_1048, n1352);
  not g2186 (n_1049, n1354);
  and g2187 (n1355, n_1048, n_1049);
  not g2188 (n_1050, n1345);
  not g2189 (n_1051, n1355);
  and g2190 (n1356, n_1050, n_1051);
  not g2191 (n_1052, n1356);
  and g2192 (n1357, n_1050, n_1052);
  and g2193 (n1358, n_1051, n_1052);
  not g2194 (n_1053, n1357);
  not g2195 (n_1054, n1358);
  and g2196 (n1359, n_1053, n_1054);
  and g2197 (n1360, n_1003, n_1007);
  and g2198 (n1361, n1359, n1360);
  not g2199 (n_1055, n1359);
  not g2200 (n_1056, n1360);
  and g2201 (n1362, n_1055, n_1056);
  not g2202 (n_1057, n1361);
  not g2203 (n_1058, n1362);
  and g2204 (n1363, n_1057, n_1058);
  and g2205 (n1364, \a[0] , \a[23] );
  and g2206 (n1365, \a[2] , \a[21] );
  not g2207 (n_1060, n1364);
  not g2208 (n_1061, n1365);
  and g2209 (n1366, n_1060, n_1061);
  and g2210 (n1367, \a[21] , \a[23] );
  and g2211 (n1368, n196, n1367);
  not g2212 (n_1062, n1366);
  not g2213 (n_1063, n1368);
  and g2214 (n1369, n_1062, n_1063);
  and g2215 (n1370, n1297, n1369);
  not g2216 (n_1064, n1370);
  and g2217 (n1371, n_1063, n_1064);
  and g2218 (n1372, n_1062, n1371);
  and g2219 (n1373, n1297, n_1064);
  not g2220 (n_1065, n1372);
  not g2221 (n_1066, n1373);
  and g2222 (n1374, n_1065, n_1066);
  not g2223 (n_1067, n1374);
  and g2224 (n1375, n1255, n_1067);
  not g2225 (n_1068, n1255);
  and g2226 (n1376, n_1068, n1374);
  not g2227 (n_1069, n1375);
  not g2228 (n_1070, n1376);
  and g2229 (n1377, n_1069, n_1070);
  and g2230 (n1378, n432, n895);
  and g2231 (n1379, n763, n893);
  and g2232 (n1380, n380, n891);
  not g2233 (n_1071, n1379);
  not g2234 (n_1072, n1380);
  and g2235 (n1381, n_1071, n_1072);
  not g2236 (n_1073, n1378);
  not g2237 (n_1074, n1381);
  and g2238 (n1382, n_1073, n_1074);
  not g2239 (n_1075, n1382);
  and g2240 (n1383, \a[16] , n_1075);
  and g2241 (n1384, \a[7] , n1383);
  and g2242 (n1385, \a[9] , \a[14] );
  not g2243 (n_1076, n1107);
  not g2244 (n_1077, n1385);
  and g2245 (n1386, n_1076, n_1077);
  and g2246 (n1387, n_1073, n_1075);
  not g2247 (n_1078, n1386);
  and g2248 (n1388, n_1078, n1387);
  not g2249 (n_1079, n1384);
  not g2250 (n_1080, n1388);
  and g2251 (n1389, n_1079, n_1080);
  not g2252 (n_1081, n1377);
  not g2253 (n_1082, n1389);
  and g2254 (n1390, n_1081, n_1082);
  and g2255 (n1391, n1377, n1389);
  not g2256 (n_1083, n1390);
  not g2257 (n_1084, n1391);
  and g2258 (n1392, n_1083, n_1084);
  not g2259 (n_1085, n1363);
  not g2260 (n_1086, n1392);
  and g2261 (n1393, n_1085, n_1086);
  and g2262 (n1394, n1363, n1392);
  not g2263 (n_1087, n1393);
  not g2264 (n_1088, n1394);
  and g2265 (n1395, n_1087, n_1088);
  not g2266 (n_1089, n1330);
  and g2267 (n1396, n_1089, n1395);
  not g2268 (n_1090, n1395);
  and g2269 (n1397, n1330, n_1090);
  not g2270 (n_1091, n1396);
  not g2271 (n_1092, n1397);
  and g2272 (n1398, n_1091, n_1092);
  and g2273 (n1399, n_958, n_997);
  and g2274 (n1400, n_949, n_954);
  and g2275 (n1401, n_976, n_991);
  and g2276 (n1402, n1400, n1401);
  not g2277 (n_1093, n1400);
  not g2278 (n_1094, n1401);
  and g2279 (n1403, n_1093, n_1094);
  not g2280 (n_1095, n1402);
  not g2281 (n_1096, n1403);
  and g2282 (n1404, n_1095, n_1096);
  and g2283 (n1405, \a[1] , \a[22] );
  and g2284 (n1406, \a[12] , n1405);
  not g2285 (n_1097, n1405);
  and g2286 (n1407, n_325, n_1097);
  not g2287 (n_1098, n1406);
  not g2288 (n_1099, n1407);
  and g2289 (n1408, n_1098, n_1099);
  not g2290 (n_1100, n1408);
  and g2291 (n1409, n1281, n_1100);
  not g2292 (n_1101, n1281);
  and g2293 (n1410, n_1101, n1408);
  not g2294 (n_1102, n1409);
  not g2295 (n_1103, n1410);
  and g2296 (n1411, n_1102, n_1103);
  not g2297 (n_1104, n1266);
  and g2298 (n1412, n_1104, n1411);
  not g2299 (n_1105, n1411);
  and g2300 (n1413, n1266, n_1105);
  not g2301 (n_1106, n1412);
  not g2302 (n_1107, n1413);
  and g2303 (n1414, n_1106, n_1107);
  and g2304 (n1415, n1404, n1414);
  not g2305 (n_1108, n1404);
  not g2306 (n_1109, n1414);
  and g2307 (n1416, n_1108, n_1109);
  not g2308 (n_1110, n1415);
  not g2309 (n_1111, n1416);
  and g2310 (n1417, n_1110, n_1111);
  not g2311 (n_1112, n1399);
  and g2312 (n1418, n_1112, n1417);
  not g2313 (n_1113, n1417);
  and g2314 (n1419, n1399, n_1113);
  not g2315 (n_1114, n1418);
  not g2316 (n_1115, n1419);
  and g2317 (n1420, n_1114, n_1115);
  and g2318 (n1421, n1398, n1420);
  not g2319 (n_1116, n1398);
  not g2320 (n_1117, n1420);
  and g2321 (n1422, n_1116, n_1117);
  not g2322 (n_1118, n1421);
  not g2323 (n_1119, n1422);
  and g2324 (n1423, n_1118, n_1119);
  not g2325 (n_1120, n1423);
  and g2326 (n1424, n1329, n_1120);
  not g2327 (n_1121, n1329);
  and g2328 (n1425, n_1121, n1423);
  not g2329 (n_1122, n1424);
  not g2330 (n_1123, n1425);
  and g2331 (n1426, n_1122, n_1123);
  not g2332 (n_1124, n1326);
  and g2333 (n1427, n_1027, n_1124);
  not g2334 (n_1125, n1426);
  and g2335 (n1428, n_1125, n1427);
  not g2336 (n_1126, n1427);
  and g2337 (n1429, n1426, n_1126);
  not g2338 (n_1127, n1428);
  not g2339 (n_1128, n1429);
  and g2340 (\asquared[24] , n_1127, n_1128);
  and g2341 (n1431, n_1122, n_1126);
  not g2342 (n_1129, n1431);
  and g2343 (n1432, n_1123, n_1129);
  and g2344 (n1433, n_1114, n_1118);
  and g2345 (n1434, n_1088, n_1091);
  and g2346 (n1435, n1338, n1353);
  not g2347 (n_1130, n1338);
  not g2348 (n_1131, n1353);
  and g2349 (n1436, n_1130, n_1131);
  not g2350 (n_1132, n1435);
  not g2351 (n_1133, n1436);
  and g2352 (n1437, n_1132, n_1133);
  not g2353 (n_1134, n1437);
  and g2354 (n1438, n1387, n_1134);
  not g2355 (n_1135, n1387);
  and g2356 (n1439, n_1135, n1437);
  not g2357 (n_1136, n1438);
  not g2358 (n_1137, n1439);
  and g2359 (n1440, n_1136, n_1137);
  and g2360 (n1441, n_1052, n_1058);
  and g2361 (n1442, n_1068, n_1067);
  not g2362 (n_1138, n1442);
  and g2363 (n1443, n_1083, n_1138);
  and g2364 (n1444, n1441, n1443);
  not g2365 (n_1139, n1441);
  not g2366 (n_1140, n1443);
  and g2367 (n1445, n_1139, n_1140);
  not g2368 (n_1141, n1444);
  not g2369 (n_1142, n1445);
  and g2370 (n1446, n_1141, n_1142);
  and g2371 (n1447, n1440, n1446);
  not g2372 (n_1143, n1440);
  not g2373 (n_1144, n1446);
  and g2374 (n1448, n_1143, n_1144);
  not g2375 (n_1145, n1447);
  not g2376 (n_1146, n1448);
  and g2377 (n1449, n_1145, n_1146);
  not g2378 (n_1147, n1434);
  and g2379 (n1450, n_1147, n1449);
  not g2380 (n_1148, n1450);
  and g2381 (n1451, n_1147, n_1148);
  and g2382 (n1452, n1449, n_1148);
  not g2383 (n_1149, n1451);
  not g2384 (n_1150, n1452);
  and g2385 (n1453, n_1149, n_1150);
  and g2386 (n1454, \a[0] , \a[24] );
  and g2387 (n1455, n1406, n1454);
  not g2388 (n_1152, n1455);
  and g2389 (n1456, n1406, n_1152);
  and g2390 (n1457, n_1098, n1454);
  not g2391 (n_1153, n1456);
  not g2392 (n_1154, n1457);
  and g2393 (n1458, n_1153, n_1154);
  and g2394 (n1459, \a[1] , \a[23] );
  and g2395 (n1460, n818, n1459);
  not g2396 (n_1155, n1460);
  and g2397 (n1461, n1459, n_1155);
  and g2398 (n1462, n818, n_1155);
  not g2399 (n_1156, n1461);
  not g2400 (n_1157, n1462);
  and g2401 (n1463, n_1156, n_1157);
  not g2402 (n_1158, n1458);
  not g2403 (n_1159, n1463);
  and g2404 (n1464, n_1158, n_1159);
  not g2405 (n_1160, n1464);
  and g2406 (n1465, n_1158, n_1160);
  and g2407 (n1466, n_1159, n_1160);
  not g2408 (n_1161, n1465);
  not g2409 (n_1162, n1466);
  and g2410 (n1467, n_1161, n_1162);
  and g2411 (n1468, \a[7] , \a[17] );
  and g2412 (n1469, \a[18] , \a[22] );
  and g2413 (n1470, n310, n1469);
  and g2414 (n1471, n335, n1052);
  and g2415 (n1472, \a[2] , \a[22] );
  and g2416 (n1473, n1468, n1472);
  not g2417 (n_1163, n1471);
  not g2418 (n_1164, n1473);
  and g2419 (n1474, n_1163, n_1164);
  not g2420 (n_1165, n1470);
  not g2421 (n_1166, n1474);
  and g2422 (n1475, n_1165, n_1166);
  not g2423 (n_1167, n1475);
  and g2424 (n1476, n1468, n_1167);
  and g2425 (n1477, n_1165, n_1167);
  and g2426 (n1478, \a[6] , \a[18] );
  not g2427 (n_1168, n1472);
  not g2428 (n_1169, n1478);
  and g2429 (n1479, n_1168, n_1169);
  not g2430 (n_1170, n1479);
  and g2431 (n1480, n1477, n_1170);
  not g2432 (n_1171, n1476);
  not g2433 (n_1172, n1480);
  and g2434 (n1481, n_1171, n_1172);
  not g2435 (n_1173, n1467);
  not g2436 (n_1174, n1481);
  and g2437 (n1482, n_1173, n_1174);
  not g2438 (n_1175, n1482);
  and g2439 (n1483, n_1173, n_1175);
  and g2440 (n1484, n_1174, n_1175);
  not g2441 (n_1176, n1483);
  not g2442 (n_1177, n1484);
  and g2443 (n1485, n_1176, n_1177);
  and g2444 (n1486, n_1103, n_1106);
  and g2445 (n1487, n1485, n1486);
  not g2446 (n_1178, n1485);
  not g2447 (n_1179, n1486);
  and g2448 (n1488, n_1178, n_1179);
  not g2449 (n_1180, n1487);
  not g2450 (n_1181, n1488);
  and g2451 (n1489, n_1180, n_1181);
  and g2452 (n1490, \a[19] , \a[20] );
  and g2453 (n1491, n226, n1490);
  and g2454 (n1492, \a[19] , \a[21] );
  and g2455 (n1493, n300, n1492);
  and g2456 (n1494, \a[20] , \a[21] );
  and g2457 (n1495, n209, n1494);
  not g2458 (n_1182, n1493);
  not g2459 (n_1183, n1495);
  and g2460 (n1496, n_1182, n_1183);
  not g2461 (n_1184, n1491);
  not g2462 (n_1185, n1496);
  and g2463 (n1497, n_1184, n_1185);
  not g2464 (n_1186, n1497);
  and g2465 (n1498, \a[3] , n_1186);
  and g2466 (n1499, \a[21] , n1498);
  and g2467 (n1500, n_1184, n_1186);
  and g2468 (n1501, \a[4] , \a[20] );
  and g2469 (n1502, \a[5] , \a[19] );
  not g2470 (n_1187, n1501);
  not g2471 (n_1188, n1502);
  and g2472 (n1503, n_1187, n_1188);
  not g2473 (n_1189, n1503);
  and g2474 (n1504, n1500, n_1189);
  not g2475 (n_1190, n1499);
  not g2476 (n_1191, n1504);
  and g2477 (n1505, n_1190, n_1191);
  not g2478 (n_1192, n1505);
  and g2479 (n1506, n1371, n_1192);
  not g2480 (n_1193, n1371);
  and g2481 (n1507, n_1193, n1505);
  not g2482 (n_1194, n1506);
  not g2483 (n_1195, n1507);
  and g2484 (n1508, n_1194, n_1195);
  and g2485 (n1509, \a[8] , \a[16] );
  and g2486 (n1510, n484, n895);
  and g2487 (n1511, n378, n893);
  and g2488 (n1512, n432, n891);
  not g2489 (n_1196, n1511);
  not g2490 (n_1197, n1512);
  and g2491 (n1513, n_1196, n_1197);
  not g2492 (n_1198, n1510);
  not g2493 (n_1199, n1513);
  and g2494 (n1514, n_1198, n_1199);
  not g2495 (n_1200, n1514);
  and g2496 (n1515, n1509, n_1200);
  and g2497 (n1516, n_1198, n_1200);
  and g2498 (n1517, \a[9] , \a[15] );
  and g2499 (n1518, \a[10] , \a[14] );
  not g2500 (n_1201, n1517);
  not g2501 (n_1202, n1518);
  and g2502 (n1519, n_1201, n_1202);
  not g2503 (n_1203, n1519);
  and g2504 (n1520, n1516, n_1203);
  not g2505 (n_1204, n1515);
  not g2506 (n_1205, n1520);
  and g2507 (n1521, n_1204, n_1205);
  not g2508 (n_1206, n1508);
  not g2509 (n_1207, n1521);
  and g2510 (n1522, n_1206, n_1207);
  and g2511 (n1523, n1508, n1521);
  not g2512 (n_1208, n1522);
  not g2513 (n_1209, n1523);
  and g2514 (n1524, n_1208, n_1209);
  not g2515 (n_1210, n1489);
  not g2516 (n_1211, n1524);
  and g2517 (n1525, n_1210, n_1211);
  and g2518 (n1526, n1489, n1524);
  not g2519 (n_1212, n1525);
  not g2520 (n_1213, n1526);
  and g2521 (n1527, n_1212, n_1213);
  and g2522 (n1528, n_1096, n_1110);
  not g2523 (n_1214, n1528);
  and g2524 (n1529, n1527, n_1214);
  not g2525 (n_1215, n1527);
  and g2526 (n1530, n_1215, n1528);
  not g2527 (n_1216, n1529);
  not g2528 (n_1217, n1530);
  and g2529 (n1531, n_1216, n_1217);
  not g2530 (n_1218, n1453);
  and g2531 (n1532, n_1218, n1531);
  not g2532 (n_1219, n1531);
  and g2533 (n1533, n_1150, n_1219);
  and g2534 (n1534, n_1149, n1533);
  not g2535 (n_1220, n1532);
  not g2536 (n_1221, n1534);
  and g2537 (n1535, n_1220, n_1221);
  not g2538 (n_1222, n1433);
  and g2539 (n1536, n_1222, n1535);
  not g2540 (n_1223, n1535);
  and g2541 (n1537, n1433, n_1223);
  not g2542 (n_1224, n1536);
  not g2543 (n_1225, n1537);
  and g2544 (n1538, n_1224, n_1225);
  not g2545 (n_1226, n1538);
  and g2546 (n1539, n1432, n_1226);
  not g2547 (n_1227, n1432);
  and g2548 (n1540, n_1227, n_1225);
  and g2549 (n1541, n_1224, n1540);
  not g2550 (n_1228, n1539);
  not g2551 (n_1229, n1541);
  and g2552 (\asquared[25] , n_1228, n_1229);
  and g2553 (n1543, n_1148, n_1220);
  and g2554 (n1544, \a[0] , \a[25] );
  and g2555 (n1545, \a[2] , \a[23] );
  not g2556 (n_1231, n1544);
  not g2557 (n_1232, n1545);
  and g2558 (n1546, n_1231, n_1232);
  and g2559 (n1547, \a[23] , \a[25] );
  and g2560 (n1548, n196, n1547);
  not g2561 (n_1233, n1548);
  and g2562 (n1549, n685, n_1233);
  not g2563 (n_1234, n1546);
  and g2564 (n1550, n_1234, n1549);
  not g2565 (n_1235, n1550);
  and g2566 (n1551, n_1233, n_1235);
  and g2567 (n1552, n_1234, n1551);
  and g2568 (n1553, n685, n_1235);
  not g2569 (n_1236, n1552);
  not g2570 (n_1237, n1553);
  and g2571 (n1554, n_1236, n_1237);
  and g2572 (n1555, n432, n1048);
  and g2573 (n1556, n763, n1050);
  and g2574 (n1557, n380, n1052);
  not g2575 (n_1238, n1556);
  not g2576 (n_1239, n1557);
  and g2577 (n1558, n_1238, n_1239);
  not g2578 (n_1240, n1555);
  not g2579 (n_1241, n1558);
  and g2580 (n1559, n_1240, n_1241);
  not g2581 (n_1242, n1559);
  and g2582 (n1560, n876, n_1242);
  and g2583 (n1561, n_1240, n_1242);
  and g2584 (n1562, \a[8] , \a[17] );
  not g2585 (n_1243, n847);
  not g2586 (n_1244, n1562);
  and g2587 (n1563, n_1243, n_1244);
  not g2588 (n_1245, n1563);
  and g2589 (n1564, n1561, n_1245);
  not g2590 (n_1246, n1560);
  not g2591 (n_1247, n1564);
  and g2592 (n1565, n_1246, n_1247);
  not g2593 (n_1248, n1554);
  not g2594 (n_1249, n1565);
  and g2595 (n1566, n_1248, n_1249);
  not g2596 (n_1250, n1566);
  and g2597 (n1567, n_1248, n_1250);
  and g2598 (n1568, n_1249, n_1250);
  not g2599 (n_1251, n1567);
  not g2600 (n_1252, n1568);
  and g2601 (n1569, n_1251, n_1252);
  and g2602 (n1570, \a[6] , \a[19] );
  and g2603 (n1571, \a[22] , n1273);
  and g2604 (n1572, \a[4] , n1492);
  not g2605 (n_1253, n1571);
  not g2606 (n_1254, n1572);
  and g2607 (n1573, n_1253, n_1254);
  and g2608 (n1574, \a[21] , \a[22] );
  and g2609 (n1575, n209, n1574);
  not g2610 (n_1255, n1575);
  and g2611 (n1576, \a[6] , n_1255);
  not g2612 (n_1256, n1573);
  and g2613 (n1577, n_1256, n1576);
  not g2614 (n_1257, n1577);
  and g2615 (n1578, n1570, n_1257);
  and g2616 (n1579, n_1255, n_1257);
  and g2617 (n1580, \a[3] , \a[22] );
  and g2618 (n1581, \a[4] , \a[21] );
  not g2619 (n_1258, n1580);
  not g2620 (n_1259, n1581);
  and g2621 (n1582, n_1258, n_1259);
  not g2622 (n_1260, n1582);
  and g2623 (n1583, n1579, n_1260);
  not g2624 (n_1261, n1578);
  not g2625 (n_1262, n1583);
  and g2626 (n1584, n_1261, n_1262);
  not g2627 (n_1263, n1569);
  not g2628 (n_1264, n1584);
  and g2629 (n1585, n_1263, n_1264);
  not g2630 (n_1265, n1585);
  and g2631 (n1586, n_1263, n_1265);
  and g2632 (n1587, n_1264, n_1265);
  not g2633 (n_1266, n1586);
  not g2634 (n_1267, n1587);
  and g2635 (n1588, n_1266, n_1267);
  and g2636 (n1589, n_1142, n_1145);
  not g2637 (n_1268, n1588);
  not g2638 (n_1269, n1589);
  and g2639 (n1590, n_1268, n_1269);
  not g2640 (n_1270, n1590);
  and g2641 (n1591, n_1268, n_1270);
  and g2642 (n1592, n_1269, n_1270);
  not g2643 (n_1271, n1591);
  not g2644 (n_1272, n1592);
  and g2645 (n1593, n_1271, n_1272);
  and g2646 (n1594, \a[1] , \a[24] );
  and g2647 (n1595, \a[13] , n1594);
  not g2648 (n_1273, \a[13] );
  not g2649 (n_1274, n1594);
  and g2650 (n1596, n_1273, n_1274);
  not g2651 (n_1275, n1595);
  not g2652 (n_1276, n1596);
  and g2653 (n1597, n_1275, n_1276);
  and g2654 (n1598, n1460, n1597);
  not g2655 (n_1277, n1597);
  and g2656 (n1599, n_1155, n_1277);
  not g2657 (n_1278, n1598);
  not g2658 (n_1279, n1599);
  and g2659 (n1600, n_1278, n_1279);
  not g2660 (n_1280, n1500);
  and g2661 (n1601, n_1280, n1600);
  not g2662 (n_1281, n1600);
  and g2663 (n1602, n1500, n_1281);
  not g2664 (n_1282, n1601);
  not g2665 (n_1283, n1602);
  and g2666 (n1603, n_1282, n_1283);
  and g2667 (n1604, n_1133, n_1137);
  and g2668 (n1605, \a[11] , \a[14] );
  not g2669 (n_1284, n748);
  not g2670 (n_1285, n1605);
  and g2671 (n1606, n_1284, n_1285);
  and g2672 (n1607, n748, n1605);
  not g2673 (n_1286, n1607);
  not g2676 (n_1287, n1606);
  not g2678 (n_1288, n1610);
  and g2679 (n1611, \a[5] , n_1288);
  and g2680 (n1612, \a[20] , n1611);
  and g2681 (n1613, n_1286, n_1288);
  and g2682 (n1614, n_1287, n1613);
  not g2683 (n_1289, n1612);
  not g2684 (n_1290, n1614);
  and g2685 (n1615, n_1289, n_1290);
  not g2686 (n_1291, n1604);
  not g2687 (n_1292, n1615);
  and g2688 (n1616, n_1291, n_1292);
  not g2689 (n_1293, n1616);
  and g2690 (n1617, n_1291, n_1293);
  and g2691 (n1618, n_1292, n_1293);
  not g2692 (n_1294, n1617);
  not g2693 (n_1295, n1618);
  and g2694 (n1619, n_1294, n_1295);
  not g2695 (n_1296, n1619);
  and g2696 (n1620, n1603, n_1296);
  not g2697 (n_1297, n1620);
  and g2698 (n1621, n1603, n_1297);
  and g2699 (n1622, n_1296, n_1297);
  not g2700 (n_1298, n1621);
  not g2701 (n_1299, n1622);
  and g2702 (n1623, n_1298, n_1299);
  not g2703 (n_1300, n1593);
  not g2704 (n_1301, n1623);
  and g2705 (n1624, n_1300, n_1301);
  not g2706 (n_1302, n1624);
  and g2707 (n1625, n_1300, n_1302);
  and g2708 (n1626, n_1301, n_1302);
  not g2709 (n_1303, n1625);
  not g2710 (n_1304, n1626);
  and g2711 (n1627, n_1303, n_1304);
  and g2712 (n1628, n1477, n1516);
  not g2713 (n_1305, n1477);
  not g2714 (n_1306, n1516);
  and g2715 (n1629, n_1305, n_1306);
  not g2716 (n_1307, n1628);
  not g2717 (n_1308, n1629);
  and g2718 (n1630, n_1307, n_1308);
  and g2719 (n1631, n_1152, n_1160);
  not g2720 (n_1309, n1630);
  and g2721 (n1632, n_1309, n1631);
  not g2722 (n_1310, n1631);
  and g2723 (n1633, n1630, n_1310);
  not g2724 (n_1311, n1632);
  not g2725 (n_1312, n1633);
  and g2726 (n1634, n_1311, n_1312);
  and g2727 (n1635, n_1193, n_1192);
  not g2728 (n_1313, n1635);
  and g2729 (n1636, n_1208, n_1313);
  not g2730 (n_1314, n1634);
  and g2731 (n1637, n_1314, n1636);
  not g2732 (n_1315, n1636);
  and g2733 (n1638, n1634, n_1315);
  not g2734 (n_1316, n1637);
  not g2735 (n_1317, n1638);
  and g2736 (n1639, n_1316, n_1317);
  and g2737 (n1640, n_1175, n_1181);
  not g2738 (n_1318, n1639);
  and g2739 (n1641, n_1318, n1640);
  not g2740 (n_1319, n1640);
  and g2741 (n1642, n1639, n_1319);
  not g2742 (n_1320, n1641);
  not g2743 (n_1321, n1642);
  and g2744 (n1643, n_1320, n_1321);
  and g2745 (n1644, n_1213, n_1216);
  not g2746 (n_1322, n1644);
  and g2747 (n1645, n1643, n_1322);
  not g2748 (n_1323, n1645);
  and g2749 (n1646, n1643, n_1323);
  and g2750 (n1647, n_1322, n_1323);
  not g2751 (n_1324, n1646);
  not g2752 (n_1325, n1647);
  and g2753 (n1648, n_1324, n_1325);
  not g2754 (n_1326, n1627);
  not g2755 (n_1327, n1648);
  and g2756 (n1649, n_1326, n_1327);
  and g2757 (n1650, n1627, n_1325);
  and g2758 (n1651, n_1324, n1650);
  not g2759 (n_1328, n1649);
  not g2760 (n_1329, n1651);
  and g2761 (n1652, n_1328, n_1329);
  not g2762 (n_1330, n1652);
  and g2763 (n1653, n1543, n_1330);
  not g2764 (n_1331, n1543);
  and g2765 (n1654, n_1331, n1652);
  not g2766 (n_1332, n1653);
  not g2767 (n_1333, n1654);
  and g2768 (n1655, n_1332, n_1333);
  not g2769 (n_1334, n1540);
  and g2770 (n1656, n_1224, n_1334);
  not g2771 (n_1335, n1655);
  and g2772 (n1657, n_1335, n1656);
  not g2773 (n_1336, n1656);
  and g2774 (n1658, n1655, n_1336);
  not g2775 (n_1337, n1657);
  not g2776 (n_1338, n1658);
  and g2777 (\asquared[26] , n_1337, n_1338);
  and g2778 (n1660, n_1323, n_1328);
  and g2779 (n1661, \a[3] , \a[23] );
  and g2780 (n1662, \a[7] , \a[19] );
  not g2781 (n_1339, n1661);
  not g2782 (n_1340, n1662);
  and g2783 (n1663, n_1339, n_1340);
  and g2784 (n1664, \a[19] , \a[24] );
  and g2785 (n1665, n343, n1664);
  and g2786 (n1666, \a[23] , \a[24] );
  and g2787 (n1667, n218, n1666);
  not g2788 (n_1341, n1665);
  not g2789 (n_1342, n1667);
  and g2790 (n1668, n_1341, n_1342);
  and g2791 (n1669, n1661, n1662);
  not g2792 (n_1343, n1668);
  not g2793 (n_1344, n1669);
  and g2794 (n1670, n_1343, n_1344);
  not g2795 (n_1345, n1670);
  and g2796 (n1671, n_1344, n_1345);
  not g2797 (n_1346, n1663);
  and g2798 (n1672, n_1346, n1671);
  and g2799 (n1673, \a[24] , n_1345);
  and g2800 (n1674, \a[2] , n1673);
  not g2801 (n_1347, n1672);
  not g2802 (n_1348, n1674);
  and g2803 (n1675, n_1347, n_1348);
  and g2804 (n1676, \a[9] , \a[17] );
  and g2805 (n1677, n723, n891);
  and g2806 (n1678, n816, n1676);
  and g2807 (n1679, n484, n1048);
  not g2808 (n_1349, n1678);
  not g2809 (n_1350, n1679);
  and g2810 (n1680, n_1349, n_1350);
  not g2811 (n_1351, n1677);
  not g2812 (n_1352, n1680);
  and g2813 (n1681, n_1351, n_1352);
  not g2814 (n_1353, n1681);
  and g2815 (n1682, n1676, n_1353);
  and g2816 (n1683, n_1351, n_1353);
  and g2817 (n1684, \a[10] , \a[16] );
  not g2818 (n_1354, n816);
  not g2819 (n_1355, n1684);
  and g2820 (n1685, n_1354, n_1355);
  not g2821 (n_1356, n1685);
  and g2822 (n1686, n1683, n_1356);
  not g2823 (n_1357, n1682);
  not g2824 (n_1358, n1686);
  and g2825 (n1687, n_1357, n_1358);
  not g2826 (n_1359, n1675);
  not g2827 (n_1360, n1687);
  and g2828 (n1688, n_1359, n_1360);
  not g2829 (n_1361, n1688);
  and g2830 (n1689, n_1359, n_1361);
  and g2831 (n1690, n_1360, n_1361);
  not g2832 (n_1362, n1689);
  not g2833 (n_1363, n1690);
  and g2834 (n1691, n_1362, n_1363);
  and g2835 (n1692, n332, n1494);
  and g2836 (n1693, \a[20] , \a[22] );
  and g2837 (n1694, n400, n1693);
  and g2838 (n1695, n226, n1574);
  not g2839 (n_1364, n1694);
  not g2840 (n_1365, n1695);
  and g2841 (n1696, n_1364, n_1365);
  not g2842 (n_1366, n1692);
  not g2843 (n_1367, n1696);
  and g2844 (n1697, n_1366, n_1367);
  not g2845 (n_1368, n1697);
  and g2846 (n1698, \a[22] , n_1368);
  and g2847 (n1699, \a[4] , n1698);
  and g2848 (n1700, n_1366, n_1368);
  and g2849 (n1701, \a[5] , \a[21] );
  and g2850 (n1702, \a[6] , \a[20] );
  not g2851 (n_1369, n1701);
  not g2852 (n_1370, n1702);
  and g2853 (n1703, n_1369, n_1370);
  not g2854 (n_1371, n1703);
  and g2855 (n1704, n1700, n_1371);
  not g2856 (n_1372, n1699);
  not g2857 (n_1373, n1704);
  and g2858 (n1705, n_1372, n_1373);
  not g2859 (n_1374, n1691);
  not g2860 (n_1375, n1705);
  and g2861 (n1706, n_1374, n_1375);
  not g2862 (n_1376, n1706);
  and g2863 (n1707, n_1374, n_1376);
  and g2864 (n1708, n_1375, n_1376);
  not g2865 (n_1377, n1707);
  not g2866 (n_1378, n1708);
  and g2867 (n1709, n_1377, n_1378);
  and g2868 (n1710, n_1317, n_1321);
  and g2869 (n1711, n1709, n1710);
  not g2870 (n_1379, n1709);
  not g2871 (n_1380, n1710);
  and g2872 (n1712, n_1379, n_1380);
  not g2873 (n_1381, n1711);
  not g2874 (n_1382, n1712);
  and g2875 (n1713, n_1381, n_1382);
  and g2876 (n1714, n_1308, n_1312);
  and g2877 (n1715, n_1278, n_1282);
  and g2878 (n1716, n1714, n1715);
  not g2879 (n_1383, n1714);
  not g2880 (n_1384, n1715);
  and g2881 (n1717, n_1383, n_1384);
  not g2882 (n_1385, n1716);
  not g2883 (n_1386, n1717);
  and g2884 (n1718, n_1385, n_1386);
  and g2885 (n1719, n1551, n1561);
  not g2886 (n_1387, n1551);
  not g2887 (n_1388, n1561);
  and g2888 (n1720, n_1387, n_1388);
  not g2889 (n_1389, n1719);
  not g2890 (n_1390, n1720);
  and g2891 (n1721, n_1389, n_1390);
  and g2892 (n1722, \a[0] , \a[26] );
  and g2893 (n1723, \a[8] , \a[18] );
  not g2894 (n_1392, n1722);
  not g2895 (n_1393, n1723);
  and g2896 (n1724, n_1392, n_1393);
  and g2897 (n1725, n1722, n1723);
  not g2898 (n_1394, n1724);
  not g2899 (n_1395, n1725);
  and g2900 (n1726, n_1394, n_1395);
  and g2901 (n1727, n1595, n1726);
  not g2902 (n_1396, n1727);
  and g2903 (n1728, n1595, n_1396);
  and g2904 (n1729, n_1395, n_1396);
  and g2905 (n1730, n_1394, n1729);
  not g2906 (n_1397, n1728);
  not g2907 (n_1398, n1730);
  and g2908 (n1731, n_1397, n_1398);
  not g2909 (n_1399, n1731);
  and g2910 (n1732, n1721, n_1399);
  not g2911 (n_1400, n1732);
  and g2912 (n1733, n1721, n_1400);
  and g2913 (n1734, n_1399, n_1400);
  not g2914 (n_1401, n1733);
  not g2915 (n_1402, n1734);
  and g2916 (n1735, n_1401, n_1402);
  not g2917 (n_1403, n1735);
  and g2918 (n1736, n1718, n_1403);
  not g2919 (n_1404, n1718);
  and g2920 (n1737, n_1404, n1735);
  not g2921 (n_1405, n1737);
  and g2922 (n1738, n1713, n_1405);
  not g2923 (n_1406, n1736);
  and g2924 (n1739, n_1406, n1738);
  not g2925 (n_1407, n1739);
  and g2926 (n1740, n1713, n_1407);
  and g2927 (n1741, n_1405, n_1407);
  and g2928 (n1742, n_1406, n1741);
  not g2929 (n_1408, n1740);
  not g2930 (n_1409, n1742);
  and g2931 (n1743, n_1408, n_1409);
  and g2932 (n1744, n_1270, n_1302);
  and g2933 (n1745, n_1293, n_1297);
  and g2934 (n1746, n_1250, n_1265);
  and g2935 (n1747, \a[1] , \a[25] );
  not g2936 (n_1410, n606);
  not g2937 (n_1411, n1747);
  and g2938 (n1748, n_1410, n_1411);
  and g2939 (n1749, n606, n1747);
  not g2940 (n_1412, n1613);
  not g2941 (n_1413, n1749);
  and g2942 (n1750, n_1412, n_1413);
  not g2943 (n_1414, n1748);
  and g2944 (n1751, n_1414, n1750);
  not g2945 (n_1415, n1751);
  and g2946 (n1752, n_1412, n_1415);
  and g2947 (n1753, n_1413, n_1415);
  and g2948 (n1754, n_1414, n1753);
  not g2949 (n_1416, n1752);
  not g2950 (n_1417, n1754);
  and g2951 (n1755, n_1416, n_1417);
  not g2952 (n_1418, n1579);
  not g2953 (n_1419, n1755);
  and g2954 (n1756, n_1418, n_1419);
  and g2955 (n1757, n1579, n_1417);
  and g2956 (n1758, n_1416, n1757);
  not g2957 (n_1420, n1756);
  not g2958 (n_1421, n1758);
  and g2959 (n1759, n_1420, n_1421);
  not g2960 (n_1422, n1746);
  and g2961 (n1760, n_1422, n1759);
  not g2962 (n_1423, n1759);
  and g2963 (n1761, n1746, n_1423);
  not g2964 (n_1424, n1760);
  not g2965 (n_1425, n1761);
  and g2966 (n1762, n_1424, n_1425);
  not g2967 (n_1426, n1745);
  and g2968 (n1763, n_1426, n1762);
  not g2969 (n_1427, n1762);
  and g2970 (n1764, n1745, n_1427);
  not g2971 (n_1428, n1763);
  not g2972 (n_1429, n1764);
  and g2973 (n1765, n_1428, n_1429);
  not g2974 (n_1430, n1744);
  and g2975 (n1766, n_1430, n1765);
  not g2976 (n_1431, n1765);
  and g2977 (n1767, n1744, n_1431);
  not g2978 (n_1432, n1766);
  not g2979 (n_1433, n1767);
  and g2980 (n1768, n_1432, n_1433);
  not g2981 (n_1434, n1743);
  not g2982 (n_1435, n1768);
  and g2983 (n1769, n_1434, n_1435);
  and g2984 (n1770, n1743, n1768);
  not g2985 (n_1436, n1769);
  not g2986 (n_1437, n1770);
  and g2987 (n1771, n_1436, n_1437);
  not g2988 (n_1438, n1660);
  not g2989 (n_1439, n1771);
  and g2990 (n1772, n_1438, n_1439);
  and g2991 (n1773, n1660, n1771);
  not g2992 (n_1440, n1772);
  not g2993 (n_1441, n1773);
  and g2994 (n1774, n_1440, n_1441);
  and g2995 (n1775, n_1332, n_1336);
  not g2996 (n_1442, n1775);
  and g2997 (n1776, n_1333, n_1442);
  not g2998 (n_1443, n1774);
  and g2999 (n1777, n_1443, n1776);
  not g3000 (n_1444, n1776);
  and g3001 (n1778, n1774, n_1444);
  not g3002 (n_1445, n1777);
  not g3003 (n_1446, n1778);
  and g3004 (\asquared[27] , n_1445, n_1446);
  and g3005 (n1780, n_1434, n1768);
  not g3006 (n_1447, n1780);
  and g3007 (n1781, n_1432, n_1447);
  and g3008 (n1782, n_1382, n_1407);
  and g3009 (n1783, \a[21] , \a[24] );
  and g3010 (n1784, n340, n1783);
  and g3011 (n1785, n209, n1666);
  not g3012 (n_1448, n1784);
  not g3013 (n_1449, n1785);
  and g3014 (n1786, n_1448, n_1449);
  and g3015 (n1787, \a[4] , \a[23] );
  and g3016 (n1788, \a[6] , \a[21] );
  and g3017 (n1789, n1787, n1788);
  not g3018 (n_1450, n1786);
  not g3019 (n_1451, n1789);
  and g3020 (n1790, n_1450, n_1451);
  not g3021 (n_1452, n1790);
  and g3022 (n1791, n_1451, n_1452);
  not g3023 (n_1453, n1787);
  not g3024 (n_1454, n1788);
  and g3025 (n1792, n_1453, n_1454);
  not g3026 (n_1455, n1792);
  and g3027 (n1793, n1791, n_1455);
  and g3028 (n1794, \a[24] , n_1452);
  and g3029 (n1795, \a[3] , n1794);
  not g3030 (n_1456, n1793);
  not g3031 (n_1457, n1795);
  and g3032 (n1796, n_1456, n_1457);
  and g3033 (n1797, \a[12] , \a[15] );
  not g3034 (n_1458, n745);
  not g3035 (n_1459, n1797);
  and g3036 (n1798, n_1458, n_1459);
  and g3037 (n1799, n748, n895);
  not g3038 (n_1460, n1799);
  not g3041 (n_1461, n1798);
  not g3043 (n_1462, n1802);
  and g3044 (n1803, \a[22] , n_1462);
  and g3045 (n1804, \a[5] , n1803);
  and g3046 (n1805, n_1460, n_1462);
  and g3047 (n1806, n_1461, n1805);
  not g3048 (n_1463, n1804);
  not g3049 (n_1464, n1806);
  and g3050 (n1807, n_1463, n_1464);
  not g3051 (n_1465, n1796);
  not g3052 (n_1466, n1807);
  and g3053 (n1808, n_1465, n_1466);
  not g3054 (n_1467, n1808);
  and g3055 (n1809, n_1465, n_1467);
  and g3056 (n1810, n_1466, n_1467);
  not g3057 (n_1468, n1809);
  not g3058 (n_1469, n1810);
  and g3059 (n1811, n_1468, n_1469);
  and g3060 (n1812, \a[0] , \a[27] );
  not g3061 (n_1471, n1812);
  and g3062 (n1813, n1749, n_1471);
  and g3063 (n1814, n_1413, n1812);
  not g3064 (n_1472, n1813);
  not g3065 (n_1473, n1814);
  and g3066 (n1815, n_1472, n_1473);
  and g3067 (n1816, \a[26] , n652);
  not g3068 (n_1474, n1816);
  and g3069 (n1817, \a[14] , n_1474);
  and g3070 (n1818, \a[1] , n_1474);
  and g3071 (n1819, \a[26] , n1818);
  not g3072 (n_1475, n1817);
  not g3073 (n_1476, n1819);
  and g3074 (n1820, n_1475, n_1476);
  not g3075 (n_1477, n1815);
  not g3076 (n_1478, n1820);
  and g3077 (n1821, n_1477, n_1478);
  and g3078 (n1822, n1815, n1820);
  not g3079 (n_1479, n1821);
  not g3080 (n_1480, n1822);
  and g3081 (n1823, n_1479, n_1480);
  and g3082 (n1824, n1811, n1823);
  not g3083 (n_1481, n1811);
  not g3084 (n_1482, n1823);
  and g3085 (n1825, n_1481, n_1482);
  not g3086 (n_1483, n1824);
  not g3087 (n_1484, n1825);
  and g3088 (n1826, n_1483, n_1484);
  and g3089 (n1827, n1683, n1700);
  not g3090 (n_1485, n1683);
  not g3091 (n_1486, n1700);
  and g3092 (n1828, n_1485, n_1486);
  not g3093 (n_1487, n1827);
  not g3094 (n_1488, n1828);
  and g3095 (n1829, n_1487, n_1488);
  not g3096 (n_1489, n1829);
  and g3097 (n1830, n1671, n_1489);
  not g3098 (n_1490, n1671);
  and g3099 (n1831, n_1490, n1829);
  not g3100 (n_1491, n1830);
  not g3101 (n_1492, n1831);
  and g3102 (n1832, n_1491, n_1492);
  and g3103 (n1833, n_1386, n_1406);
  not g3104 (n_1493, n1833);
  and g3105 (n1834, n1832, n_1493);
  not g3106 (n_1494, n1832);
  and g3107 (n1835, n_1494, n1833);
  not g3108 (n_1495, n1834);
  not g3109 (n_1496, n1835);
  and g3110 (n1836, n_1495, n_1496);
  not g3111 (n_1497, n1826);
  and g3112 (n1837, n_1497, n1836);
  not g3113 (n_1498, n1836);
  and g3114 (n1838, n1826, n_1498);
  not g3115 (n_1499, n1837);
  not g3116 (n_1500, n1838);
  and g3117 (n1839, n_1499, n_1500);
  not g3118 (n_1501, n1782);
  and g3119 (n1840, n_1501, n1839);
  not g3120 (n_1502, n1839);
  and g3121 (n1841, n1782, n_1502);
  not g3122 (n_1503, n1840);
  not g3123 (n_1504, n1841);
  and g3124 (n1842, n_1503, n_1504);
  and g3125 (n1843, \a[11] , \a[16] );
  and g3126 (n1844, \a[20] , \a[25] );
  and g3127 (n1845, n343, n1844);
  and g3128 (n1846, \a[2] , \a[25] );
  and g3129 (n1847, \a[7] , \a[20] );
  not g3130 (n_1505, n1846);
  not g3131 (n_1506, n1847);
  and g3132 (n1848, n_1505, n_1506);
  not g3133 (n_1507, n1845);
  not g3134 (n_1508, n1848);
  and g3135 (n1849, n_1507, n_1508);
  not g3136 (n_1509, n1843);
  not g3137 (n_1510, n1849);
  and g3138 (n1850, n_1509, n_1510);
  and g3139 (n1851, n1843, n1849);
  not g3140 (n_1511, n1850);
  not g3141 (n_1512, n1851);
  and g3142 (n1852, n_1511, n_1512);
  not g3143 (n_1513, n1729);
  and g3144 (n1853, n_1513, n1852);
  not g3145 (n_1514, n1852);
  and g3146 (n1854, n1729, n_1514);
  not g3147 (n_1515, n1853);
  not g3148 (n_1516, n1854);
  and g3149 (n1855, n_1515, n_1516);
  and g3150 (n1856, \a[8] , \a[19] );
  and g3151 (n1857, n484, n1052);
  and g3152 (n1858, \a[10] , \a[17] );
  and g3153 (n1859, n1856, n1858);
  and g3154 (n1860, n432, n1149);
  not g3155 (n_1517, n1859);
  not g3156 (n_1518, n1860);
  and g3157 (n1861, n_1517, n_1518);
  not g3158 (n_1519, n1857);
  not g3159 (n_1520, n1861);
  and g3160 (n1862, n_1519, n_1520);
  not g3161 (n_1521, n1862);
  and g3162 (n1863, n1856, n_1521);
  and g3163 (n1864, n_1519, n_1521);
  and g3164 (n1865, \a[9] , \a[18] );
  not g3165 (n_1522, n1858);
  not g3166 (n_1523, n1865);
  and g3167 (n1866, n_1522, n_1523);
  not g3168 (n_1524, n1866);
  and g3169 (n1867, n1864, n_1524);
  not g3170 (n_1525, n1863);
  not g3171 (n_1526, n1867);
  and g3172 (n1868, n_1525, n_1526);
  not g3173 (n_1527, n1868);
  and g3174 (n1869, n1855, n_1527);
  not g3175 (n_1528, n1869);
  and g3176 (n1870, n1855, n_1528);
  and g3177 (n1871, n_1527, n_1528);
  not g3178 (n_1529, n1870);
  not g3179 (n_1530, n1871);
  and g3180 (n1872, n_1529, n_1530);
  and g3181 (n1873, n_1424, n_1428);
  and g3182 (n1874, n1872, n1873);
  not g3183 (n_1531, n1872);
  not g3184 (n_1532, n1873);
  and g3185 (n1875, n_1531, n_1532);
  not g3186 (n_1533, n1874);
  not g3187 (n_1534, n1875);
  and g3188 (n1876, n_1533, n_1534);
  and g3189 (n1877, n_1415, n_1420);
  and g3190 (n1878, n_1390, n_1400);
  and g3191 (n1879, n1877, n1878);
  not g3192 (n_1535, n1877);
  not g3193 (n_1536, n1878);
  and g3194 (n1880, n_1535, n_1536);
  not g3195 (n_1537, n1879);
  not g3196 (n_1538, n1880);
  and g3197 (n1881, n_1537, n_1538);
  and g3198 (n1882, n_1361, n_1376);
  not g3199 (n_1539, n1881);
  and g3200 (n1883, n_1539, n1882);
  not g3201 (n_1540, n1882);
  and g3202 (n1884, n1881, n_1540);
  not g3203 (n_1541, n1883);
  not g3204 (n_1542, n1884);
  and g3205 (n1885, n_1541, n_1542);
  and g3206 (n1886, n1876, n1885);
  not g3207 (n_1543, n1876);
  not g3208 (n_1544, n1885);
  and g3209 (n1887, n_1543, n_1544);
  not g3210 (n_1545, n1886);
  not g3211 (n_1546, n1887);
  and g3212 (n1888, n_1545, n_1546);
  and g3213 (n1889, n1842, n1888);
  not g3214 (n_1547, n1842);
  not g3215 (n_1548, n1888);
  and g3216 (n1890, n_1547, n_1548);
  not g3217 (n_1549, n1889);
  not g3218 (n_1550, n1890);
  and g3219 (n1891, n_1549, n_1550);
  not g3220 (n_1551, n1781);
  and g3221 (n1892, n_1551, n1891);
  not g3222 (n_1552, n1891);
  and g3223 (n1893, n1781, n_1552);
  not g3224 (n_1553, n1892);
  not g3225 (n_1554, n1893);
  and g3226 (n1894, n_1553, n_1554);
  and g3227 (n1895, n_1441, n_1444);
  not g3228 (n_1555, n1895);
  and g3229 (n1896, n_1440, n_1555);
  not g3230 (n_1556, n1894);
  and g3231 (n1897, n_1556, n1896);
  not g3232 (n_1557, n1896);
  and g3233 (n1898, n1894, n_1557);
  not g3234 (n_1558, n1897);
  not g3235 (n_1559, n1898);
  and g3236 (\asquared[28] , n_1558, n_1559);
  and g3237 (n1900, n_1495, n_1499);
  and g3238 (n1901, \a[3] , \a[25] );
  and g3239 (n1902, \a[4] , \a[24] );
  not g3240 (n_1560, n1901);
  not g3241 (n_1561, n1902);
  and g3242 (n1903, n_1560, n_1561);
  and g3243 (n1904, \a[24] , \a[25] );
  and g3244 (n1905, n209, n1904);
  not g3245 (n_1562, n1905);
  not g3248 (n_1563, n1903);
  not g3250 (n_1564, n1908);
  and g3251 (n1909, \a[8] , n_1564);
  and g3252 (n1910, \a[20] , n1909);
  and g3253 (n1911, n_1562, n_1564);
  and g3254 (n1912, n_1563, n1911);
  not g3255 (n_1565, n1910);
  not g3256 (n_1566, n1912);
  and g3257 (n1913, n_1565, n_1566);
  and g3258 (n1914, n1749, n1812);
  not g3259 (n_1567, n1914);
  and g3260 (n1915, n_1479, n_1567);
  not g3261 (n_1568, n1913);
  and g3262 (n1916, n_1568, n1915);
  not g3263 (n_1569, n1915);
  and g3264 (n1917, n1913, n_1569);
  not g3265 (n_1570, n1916);
  not g3266 (n_1571, n1917);
  and g3267 (n1918, n_1570, n_1571);
  and g3268 (n1919, \a[22] , \a[23] );
  and g3269 (n1920, n332, n1919);
  and g3270 (n1921, n268, n1367);
  and g3271 (n1922, n335, n1574);
  not g3272 (n_1572, n1921);
  not g3273 (n_1573, n1922);
  and g3274 (n1923, n_1572, n_1573);
  not g3275 (n_1574, n1920);
  not g3276 (n_1575, n1923);
  and g3277 (n1924, n_1574, n_1575);
  not g3278 (n_1576, n1924);
  and g3279 (n1925, \a[21] , n_1576);
  and g3280 (n1926, \a[7] , n1925);
  and g3281 (n1927, n_1574, n_1576);
  and g3282 (n1928, \a[5] , \a[23] );
  and g3283 (n1929, \a[6] , \a[22] );
  not g3284 (n_1577, n1928);
  not g3285 (n_1578, n1929);
  and g3286 (n1930, n_1577, n_1578);
  not g3287 (n_1579, n1930);
  and g3288 (n1931, n1927, n_1579);
  not g3289 (n_1580, n1926);
  not g3290 (n_1581, n1931);
  and g3291 (n1932, n_1580, n_1581);
  not g3292 (n_1582, n1918);
  not g3293 (n_1583, n1932);
  and g3294 (n1933, n_1582, n_1583);
  and g3295 (n1934, n1918, n1932);
  not g3296 (n_1584, n1933);
  not g3297 (n_1585, n1934);
  and g3298 (n1935, n_1584, n_1585);
  not g3299 (n_1586, n1935);
  and g3300 (n1936, n1900, n_1586);
  not g3301 (n_1587, n1900);
  and g3302 (n1937, n_1587, n1935);
  not g3303 (n_1588, n1936);
  not g3304 (n_1589, n1937);
  and g3305 (n1938, n_1588, n_1589);
  and g3306 (n1939, n_1481, n1823);
  not g3307 (n_1590, n1939);
  and g3308 (n1940, n_1467, n_1590);
  and g3309 (n1941, n_1515, n_1528);
  and g3310 (n1942, \a[1] , \a[27] );
  and g3311 (n1943, n821, n1942);
  not g3312 (n_1591, n821);
  not g3313 (n_1592, n1942);
  and g3314 (n1944, n_1591, n_1592);
  not g3315 (n_1593, n1943);
  not g3316 (n_1594, n1944);
  and g3317 (n1945, n_1593, n_1594);
  and g3318 (n1946, n1816, n1945);
  not g3319 (n_1595, n1946);
  and g3320 (n1947, n1816, n_1595);
  and g3321 (n1948, n_1474, n1945);
  not g3322 (n_1596, n1947);
  not g3323 (n_1597, n1948);
  and g3324 (n1949, n_1596, n_1597);
  not g3325 (n_1598, n1805);
  not g3326 (n_1599, n1949);
  and g3327 (n1950, n_1598, n_1599);
  and g3328 (n1951, n1805, n_1597);
  and g3329 (n1952, n_1596, n1951);
  not g3330 (n_1600, n1950);
  not g3331 (n_1601, n1952);
  and g3332 (n1953, n_1600, n_1601);
  not g3333 (n_1602, n1941);
  and g3334 (n1954, n_1602, n1953);
  not g3335 (n_1603, n1953);
  and g3336 (n1955, n1941, n_1603);
  not g3337 (n_1604, n1954);
  not g3338 (n_1605, n1955);
  and g3339 (n1956, n_1604, n_1605);
  not g3340 (n_1606, n1940);
  and g3341 (n1957, n_1606, n1956);
  not g3342 (n_1607, n1956);
  and g3343 (n1958, n1940, n_1607);
  not g3344 (n_1608, n1957);
  not g3345 (n_1609, n1958);
  and g3346 (n1959, n_1608, n_1609);
  and g3347 (n1960, n1938, n1959);
  not g3348 (n_1610, n1938);
  not g3349 (n_1611, n1959);
  and g3350 (n1961, n_1610, n_1611);
  not g3351 (n_1612, n1960);
  not g3352 (n_1613, n1961);
  and g3353 (n1962, n_1612, n_1613);
  and g3354 (n1963, n_1503, n_1549);
  and g3355 (n1964, n_1534, n_1545);
  and g3356 (n1965, n1791, n1864);
  not g3357 (n_1614, n1791);
  not g3358 (n_1615, n1864);
  and g3359 (n1966, n_1614, n_1615);
  not g3360 (n_1616, n1965);
  not g3361 (n_1617, n1966);
  and g3362 (n1967, n_1616, n_1617);
  and g3363 (n1968, n_1507, n_1512);
  not g3364 (n_1618, n1967);
  and g3365 (n1969, n_1618, n1968);
  not g3366 (n_1619, n1968);
  and g3367 (n1970, n1967, n_1619);
  not g3368 (n_1620, n1969);
  not g3369 (n_1621, n1970);
  and g3370 (n1971, n_1620, n_1621);
  and g3371 (n1972, n_1538, n_1542);
  not g3372 (n_1622, n1971);
  and g3373 (n1973, n_1622, n1972);
  not g3374 (n_1623, n1972);
  and g3375 (n1974, n1971, n_1623);
  not g3376 (n_1624, n1973);
  not g3377 (n_1625, n1974);
  and g3378 (n1975, n_1624, n_1625);
  and g3379 (n1976, \a[11] , \a[28] );
  and g3380 (n1977, n793, n1976);
  and g3381 (n1978, n602, n1048);
  not g3382 (n_1627, n1977);
  not g3383 (n_1628, n1978);
  and g3384 (n1979, n_1627, n_1628);
  and g3385 (n1980, \a[0] , \a[28] );
  and g3386 (n1981, \a[12] , \a[16] );
  and g3387 (n1982, n1980, n1981);
  not g3388 (n_1629, n1979);
  not g3389 (n_1630, n1982);
  and g3390 (n1983, n_1629, n_1630);
  not g3391 (n_1631, n1983);
  and g3392 (n1984, n_1630, n_1631);
  not g3393 (n_1632, n1980);
  not g3394 (n_1633, n1981);
  and g3395 (n1985, n_1632, n_1633);
  not g3396 (n_1634, n1985);
  and g3397 (n1986, n1984, n_1634);
  and g3398 (n1987, \a[17] , n_1631);
  and g3399 (n1988, \a[11] , n1987);
  not g3400 (n_1635, n1986);
  not g3401 (n_1636, n1988);
  and g3402 (n1989, n_1635, n_1636);
  and g3403 (n1990, \a[2] , \a[26] );
  and g3404 (n1991, \a[9] , \a[19] );
  and g3405 (n1992, \a[10] , \a[18] );
  not g3406 (n_1637, n1991);
  not g3407 (n_1638, n1992);
  and g3408 (n1993, n_1637, n_1638);
  and g3409 (n1994, n484, n1149);
  not g3410 (n_1639, n1994);
  and g3411 (n1995, n1990, n_1639);
  not g3412 (n_1640, n1993);
  and g3413 (n1996, n_1640, n1995);
  not g3414 (n_1641, n1996);
  and g3415 (n1997, n1990, n_1641);
  and g3416 (n1998, n_1639, n_1641);
  and g3417 (n1999, n_1640, n1998);
  not g3418 (n_1642, n1997);
  not g3419 (n_1643, n1999);
  and g3420 (n2000, n_1642, n_1643);
  not g3421 (n_1644, n1989);
  not g3422 (n_1645, n2000);
  and g3423 (n2001, n_1644, n_1645);
  not g3424 (n_1646, n2001);
  and g3425 (n2002, n_1644, n_1646);
  and g3426 (n2003, n_1645, n_1646);
  not g3427 (n_1647, n2002);
  not g3428 (n_1648, n2003);
  and g3429 (n2004, n_1647, n_1648);
  and g3430 (n2005, n_1488, n_1492);
  and g3431 (n2006, n2004, n2005);
  not g3432 (n_1649, n2004);
  not g3433 (n_1650, n2005);
  and g3434 (n2007, n_1649, n_1650);
  not g3435 (n_1651, n2006);
  not g3436 (n_1652, n2007);
  and g3437 (n2008, n_1651, n_1652);
  and g3438 (n2009, n1975, n2008);
  not g3439 (n_1653, n1975);
  not g3440 (n_1654, n2008);
  and g3441 (n2010, n_1653, n_1654);
  not g3442 (n_1655, n2009);
  not g3443 (n_1656, n2010);
  and g3444 (n2011, n_1655, n_1656);
  not g3445 (n_1657, n1964);
  and g3446 (n2012, n_1657, n2011);
  not g3447 (n_1658, n2011);
  and g3448 (n2013, n1964, n_1658);
  not g3449 (n_1659, n2012);
  not g3450 (n_1660, n2013);
  and g3451 (n2014, n_1659, n_1660);
  not g3452 (n_1661, n1963);
  and g3453 (n2015, n_1661, n2014);
  not g3454 (n_1662, n2014);
  and g3455 (n2016, n1963, n_1662);
  not g3456 (n_1663, n2015);
  not g3457 (n_1664, n2016);
  and g3458 (n2017, n_1663, n_1664);
  not g3459 (n_1665, n1962);
  not g3460 (n_1666, n2017);
  and g3461 (n2018, n_1665, n_1666);
  and g3462 (n2019, n1962, n2017);
  not g3463 (n_1667, n2018);
  not g3464 (n_1668, n2019);
  and g3465 (n2020, n_1667, n_1668);
  and g3466 (n2021, n_1554, n_1557);
  not g3467 (n_1669, n2021);
  and g3468 (n2022, n_1553, n_1669);
  not g3469 (n_1670, n2020);
  and g3470 (n2023, n_1670, n2022);
  not g3471 (n_1671, n2022);
  and g3472 (n2024, n2020, n_1671);
  not g3473 (n_1672, n2023);
  not g3474 (n_1673, n2024);
  and g3475 (\asquared[29] , n_1672, n_1673);
  and g3476 (n2026, n_1659, n_1663);
  and g3477 (n2027, n_1625, n_1655);
  and g3478 (n2028, n_1604, n_1608);
  and g3479 (n2029, n2027, n2028);
  not g3480 (n_1674, n2027);
  not g3481 (n_1675, n2028);
  and g3482 (n2030, n_1674, n_1675);
  not g3483 (n_1676, n2029);
  not g3484 (n_1677, n2030);
  and g3485 (n2031, n_1676, n_1677);
  and g3486 (n2032, n_1646, n_1652);
  and g3487 (n2033, n_1568, n_1569);
  not g3488 (n_1678, n2033);
  and g3489 (n2034, n_1584, n_1678);
  and g3490 (n2035, n2032, n2034);
  not g3491 (n_1679, n2032);
  not g3492 (n_1680, n2034);
  and g3493 (n2036, n_1679, n_1680);
  not g3494 (n_1681, n2035);
  not g3495 (n_1682, n2036);
  and g3496 (n2037, n_1681, n_1682);
  and g3497 (n2038, n1984, n1998);
  not g3498 (n_1683, n1984);
  not g3499 (n_1684, n1998);
  and g3500 (n2039, n_1683, n_1684);
  not g3501 (n_1685, n2038);
  not g3502 (n_1686, n2039);
  and g3503 (n2040, n_1685, n_1686);
  and g3504 (n2041, \a[27] , \a[29] );
  and g3505 (n2042, n196, n2041);
  and g3506 (n2043, \a[0] , \a[29] );
  and g3507 (n2044, \a[2] , \a[27] );
  not g3508 (n_1688, n2043);
  not g3509 (n_1689, n2044);
  and g3510 (n2045, n_1688, n_1689);
  not g3511 (n_1690, n2042);
  not g3512 (n_1691, n2045);
  and g3513 (n2046, n_1690, n_1691);
  and g3514 (n2047, n1943, n2046);
  not g3515 (n_1692, n2047);
  and g3516 (n2048, n1943, n_1692);
  and g3517 (n2049, n_1690, n_1692);
  and g3518 (n2050, n_1691, n2049);
  not g3519 (n_1693, n2048);
  not g3520 (n_1694, n2050);
  and g3521 (n2051, n_1693, n_1694);
  not g3522 (n_1695, n2051);
  and g3523 (n2052, n2040, n_1695);
  not g3524 (n_1696, n2052);
  and g3525 (n2053, n2040, n_1696);
  and g3526 (n2054, n_1695, n_1696);
  not g3527 (n_1697, n2053);
  not g3528 (n_1698, n2054);
  and g3529 (n2055, n_1697, n_1698);
  not g3530 (n_1699, n2055);
  and g3531 (n2056, n2037, n_1699);
  not g3532 (n_1700, n2037);
  and g3533 (n2057, n_1700, n2055);
  not g3534 (n_1701, n2057);
  and g3535 (n2058, n2031, n_1701);
  not g3536 (n_1702, n2056);
  and g3537 (n2059, n_1702, n2058);
  not g3538 (n_1703, n2059);
  and g3539 (n2060, n2031, n_1703);
  and g3540 (n2061, n_1701, n_1703);
  and g3541 (n2062, n_1702, n2061);
  not g3542 (n_1704, n2060);
  not g3543 (n_1705, n2062);
  and g3544 (n2063, n_1704, n_1705);
  and g3545 (n2064, n_1589, n_1612);
  and g3546 (n2065, n_1595, n_1600);
  and g3547 (n2066, \a[6] , \a[23] );
  and g3548 (n2067, \a[13] , \a[16] );
  not g3549 (n_1706, n895);
  not g3550 (n_1707, n2067);
  and g3551 (n2068, n_1706, n_1707);
  and g3552 (n2069, n895, n2067);
  not g3553 (n_1708, n2069);
  and g3554 (n2070, n2066, n_1708);
  not g3555 (n_1709, n2068);
  and g3556 (n2071, n_1709, n2070);
  not g3557 (n_1710, n2071);
  and g3558 (n2072, n2066, n_1710);
  and g3559 (n2073, n_1708, n_1710);
  and g3560 (n2074, n_1709, n2073);
  not g3561 (n_1711, n2072);
  not g3562 (n_1712, n2074);
  and g3563 (n2075, n_1711, n_1712);
  not g3564 (n_1713, n2065);
  not g3565 (n_1714, n2075);
  and g3566 (n2076, n_1713, n_1714);
  not g3567 (n_1715, n2076);
  and g3568 (n2077, n_1713, n_1715);
  and g3569 (n2078, n_1714, n_1715);
  not g3570 (n_1716, n2077);
  not g3571 (n_1717, n2078);
  and g3572 (n2079, n_1716, n_1717);
  and g3573 (n2080, n_1617, n_1621);
  and g3574 (n2081, n2079, n2080);
  not g3575 (n_1718, n2079);
  not g3576 (n_1719, n2080);
  and g3577 (n2082, n_1718, n_1719);
  not g3578 (n_1720, n2081);
  not g3579 (n_1721, n2082);
  and g3580 (n2083, n_1720, n_1721);
  and g3581 (n2084, \a[3] , \a[26] );
  and g3582 (n2085, \a[8] , \a[21] );
  not g3583 (n_1722, n2084);
  not g3584 (n_1723, n2085);
  and g3585 (n2086, n_1722, n_1723);
  and g3586 (n2087, \a[21] , \a[26] );
  and g3587 (n2088, n435, n2087);
  not g3588 (n_1724, n2088);
  not g3591 (n_1725, n2086);
  not g3593 (n_1726, n2091);
  and g3594 (n2092, n_1724, n_1726);
  and g3595 (n2093, n_1725, n2092);
  and g3596 (n2094, \a[17] , n_1726);
  and g3597 (n2095, \a[12] , n2094);
  not g3598 (n_1727, n2093);
  not g3599 (n_1728, n2095);
  and g3600 (n2096, n_1727, n_1728);
  and g3601 (n2097, n723, n1149);
  and g3602 (n2098, n1076, n1331);
  and g3603 (n2099, n484, n1490);
  not g3604 (n_1729, n2098);
  not g3605 (n_1730, n2099);
  and g3606 (n2100, n_1729, n_1730);
  not g3607 (n_1731, n2097);
  not g3608 (n_1732, n2100);
  and g3609 (n2101, n_1731, n_1732);
  not g3610 (n_1733, n2101);
  and g3611 (n2102, \a[20] , n_1733);
  and g3612 (n2103, \a[9] , n2102);
  and g3613 (n2104, n_1731, n_1733);
  and g3614 (n2105, \a[10] , \a[19] );
  and g3615 (n2106, \a[11] , \a[18] );
  not g3616 (n_1734, n2105);
  not g3617 (n_1735, n2106);
  and g3618 (n2107, n_1734, n_1735);
  not g3619 (n_1736, n2107);
  and g3620 (n2108, n2104, n_1736);
  not g3621 (n_1737, n2103);
  not g3622 (n_1738, n2108);
  and g3623 (n2109, n_1737, n_1738);
  not g3624 (n_1739, n2096);
  not g3625 (n_1740, n2109);
  and g3626 (n2110, n_1739, n_1740);
  not g3627 (n_1741, n2110);
  and g3628 (n2111, n_1739, n_1741);
  and g3629 (n2112, n_1740, n_1741);
  not g3630 (n_1742, n2111);
  not g3631 (n_1743, n2112);
  and g3632 (n2113, n_1742, n_1743);
  and g3633 (n2114, \a[4] , \a[25] );
  and g3634 (n2115, \a[22] , \a[24] );
  and g3635 (n2116, n268, n2115);
  and g3636 (n2117, n226, n1904);
  and g3637 (n2118, \a[7] , \a[22] );
  and g3638 (n2119, n2114, n2118);
  not g3639 (n_1744, n2117);
  not g3640 (n_1745, n2119);
  and g3641 (n2120, n_1744, n_1745);
  not g3642 (n_1746, n2116);
  not g3643 (n_1747, n2120);
  and g3644 (n2121, n_1746, n_1747);
  not g3645 (n_1748, n2121);
  and g3646 (n2122, n2114, n_1748);
  and g3647 (n2123, n_1746, n_1748);
  and g3648 (n2124, \a[5] , \a[24] );
  not g3649 (n_1749, n2118);
  not g3650 (n_1750, n2124);
  and g3651 (n2125, n_1749, n_1750);
  not g3652 (n_1751, n2125);
  and g3653 (n2126, n2123, n_1751);
  not g3654 (n_1752, n2122);
  not g3655 (n_1753, n2126);
  and g3656 (n2127, n_1752, n_1753);
  not g3657 (n_1754, n2113);
  not g3658 (n_1755, n2127);
  and g3659 (n2128, n_1754, n_1755);
  not g3660 (n_1756, n2128);
  and g3661 (n2129, n_1754, n_1756);
  and g3662 (n2130, n_1755, n_1756);
  not g3663 (n_1757, n2129);
  not g3664 (n_1758, n2130);
  and g3665 (n2131, n_1757, n_1758);
  and g3666 (n2132, \a[28] , n764);
  and g3667 (n2133, \a[1] , \a[28] );
  not g3668 (n_1759, \a[15] );
  not g3669 (n_1760, n2133);
  and g3670 (n2134, n_1759, n_1760);
  not g3671 (n_1761, n2132);
  not g3672 (n_1762, n2134);
  and g3673 (n2135, n_1761, n_1762);
  not g3674 (n_1763, n2135);
  and g3675 (n2136, n1927, n_1763);
  not g3676 (n_1764, n1927);
  and g3677 (n2137, n_1764, n2135);
  not g3678 (n_1765, n2136);
  not g3679 (n_1766, n2137);
  and g3680 (n2138, n_1765, n_1766);
  not g3681 (n_1767, n1911);
  and g3682 (n2139, n_1767, n2138);
  not g3683 (n_1768, n2138);
  and g3684 (n2140, n1911, n_1768);
  not g3685 (n_1769, n2139);
  not g3686 (n_1770, n2140);
  and g3687 (n2141, n_1769, n_1770);
  not g3688 (n_1771, n2131);
  and g3689 (n2142, n_1771, n2141);
  not g3690 (n_1772, n2141);
  and g3691 (n2143, n2131, n_1772);
  not g3692 (n_1773, n2142);
  not g3693 (n_1774, n2143);
  and g3694 (n2144, n_1773, n_1774);
  and g3695 (n2145, n2083, n2144);
  not g3696 (n_1775, n2083);
  not g3697 (n_1776, n2144);
  and g3698 (n2146, n_1775, n_1776);
  not g3699 (n_1777, n2145);
  not g3700 (n_1778, n2146);
  and g3701 (n2147, n_1777, n_1778);
  not g3702 (n_1779, n2064);
  and g3703 (n2148, n_1779, n2147);
  not g3704 (n_1780, n2148);
  and g3705 (n2149, n_1779, n_1780);
  and g3706 (n2150, n2147, n_1780);
  not g3707 (n_1781, n2149);
  not g3708 (n_1782, n2150);
  and g3709 (n2151, n_1781, n_1782);
  not g3710 (n_1783, n2063);
  not g3711 (n_1784, n2151);
  and g3712 (n2152, n_1783, n_1784);
  and g3713 (n2153, n2063, n_1782);
  and g3714 (n2154, n_1781, n2153);
  not g3715 (n_1785, n2152);
  not g3716 (n_1786, n2154);
  and g3717 (n2155, n_1785, n_1786);
  not g3718 (n_1787, n2026);
  and g3719 (n2156, n_1787, n2155);
  not g3720 (n_1788, n2155);
  and g3721 (n2157, n2026, n_1788);
  not g3722 (n_1789, n2156);
  not g3723 (n_1790, n2157);
  and g3724 (n2158, n_1789, n_1790);
  and g3725 (n2159, n_1667, n_1671);
  not g3726 (n_1791, n2159);
  and g3727 (n2160, n_1668, n_1791);
  not g3728 (n_1792, n2158);
  and g3729 (n2161, n_1792, n2160);
  not g3730 (n_1793, n2160);
  and g3731 (n2162, n2158, n_1793);
  not g3732 (n_1794, n2161);
  not g3733 (n_1795, n2162);
  and g3734 (\asquared[30] , n_1794, n_1795);
  and g3735 (n2164, n_1780, n_1785);
  and g3736 (n2165, \a[0] , \a[30] );
  and g3737 (n2166, n2132, n2165);
  not g3738 (n_1797, n2166);
  and g3739 (n2167, n2132, n_1797);
  and g3740 (n2168, n_1761, n2165);
  not g3741 (n_1798, n2167);
  not g3742 (n_1799, n2168);
  and g3743 (n2169, n_1798, n_1799);
  and g3744 (n2170, \a[1] , \a[29] );
  and g3745 (n2171, n893, n2170);
  not g3746 (n_1800, n2171);
  and g3747 (n2172, n2170, n_1800);
  and g3748 (n2173, n893, n_1800);
  not g3749 (n_1801, n2172);
  not g3750 (n_1802, n2173);
  and g3751 (n2174, n_1801, n_1802);
  not g3752 (n_1803, n2169);
  not g3753 (n_1804, n2174);
  and g3754 (n2175, n_1803, n_1804);
  not g3755 (n_1805, n2175);
  and g3756 (n2176, n_1803, n_1805);
  and g3757 (n2177, n_1804, n_1805);
  not g3758 (n_1806, n2176);
  not g3759 (n_1807, n2177);
  and g3760 (n2178, n_1806, n_1807);
  and g3761 (n2179, n_1766, n_1769);
  and g3762 (n2180, n2178, n2179);
  not g3763 (n_1808, n2178);
  not g3764 (n_1809, n2179);
  and g3765 (n2181, n_1808, n_1809);
  not g3766 (n_1810, n2180);
  not g3767 (n_1811, n2181);
  and g3768 (n2182, n_1810, n_1811);
  and g3769 (n2183, n_1686, n_1696);
  not g3770 (n_1812, n2182);
  and g3771 (n2184, n_1812, n2183);
  not g3772 (n_1813, n2183);
  and g3773 (n2185, n2182, n_1813);
  not g3774 (n_1814, n2184);
  not g3775 (n_1815, n2185);
  and g3776 (n2186, n_1814, n_1815);
  and g3777 (n2187, n_1773, n_1777);
  not g3778 (n_1816, n2186);
  and g3779 (n2188, n_1816, n2187);
  not g3780 (n_1817, n2187);
  and g3781 (n2189, n2186, n_1817);
  not g3782 (n_1818, n2188);
  not g3783 (n_1819, n2189);
  and g3784 (n2190, n_1818, n_1819);
  and g3785 (n2191, n2073, n2123);
  not g3786 (n_1820, n2073);
  not g3787 (n_1821, n2123);
  and g3788 (n2192, n_1820, n_1821);
  not g3789 (n_1822, n2191);
  not g3790 (n_1823, n2192);
  and g3791 (n2193, n_1822, n_1823);
  and g3792 (n2194, \a[2] , \a[28] );
  and g3793 (n2195, \a[9] , \a[21] );
  not g3794 (n_1824, n2194);
  not g3795 (n_1825, n2195);
  and g3796 (n2196, n_1824, n_1825);
  and g3797 (n2197, n2194, n2195);
  not g3798 (n_1826, n2197);
  not g3801 (n_1827, n2196);
  not g3803 (n_1828, n2200);
  and g3804 (n2201, \a[17] , n_1828);
  and g3805 (n2202, \a[13] , n2201);
  and g3806 (n2203, n_1826, n_1828);
  and g3807 (n2204, n_1827, n2203);
  not g3808 (n_1829, n2202);
  not g3809 (n_1830, n2204);
  and g3810 (n2205, n_1829, n_1830);
  not g3811 (n_1831, n2205);
  and g3812 (n2206, n2193, n_1831);
  not g3813 (n_1832, n2206);
  and g3814 (n2207, n2193, n_1832);
  and g3815 (n2208, n_1831, n_1832);
  not g3816 (n_1833, n2207);
  not g3817 (n_1834, n2208);
  and g3818 (n2209, n_1833, n_1834);
  and g3819 (n2210, n_1741, n_1756);
  and g3820 (n2211, n2209, n2210);
  not g3821 (n_1835, n2209);
  not g3822 (n_1836, n2210);
  and g3823 (n2212, n_1835, n_1836);
  not g3824 (n_1837, n2211);
  not g3825 (n_1838, n2212);
  and g3826 (n2213, n_1837, n_1838);
  and g3827 (n2214, n2092, n2104);
  not g3828 (n_1839, n2092);
  not g3829 (n_1840, n2104);
  and g3830 (n2215, n_1839, n_1840);
  not g3831 (n_1841, n2214);
  not g3832 (n_1842, n2215);
  and g3833 (n2216, n_1841, n_1842);
  not g3834 (n_1843, n2216);
  and g3835 (n2217, n2049, n_1843);
  not g3836 (n_1844, n2049);
  and g3837 (n2218, n_1844, n2216);
  not g3838 (n_1845, n2217);
  not g3839 (n_1846, n2218);
  and g3840 (n2219, n_1845, n_1846);
  and g3841 (n2220, n2213, n2219);
  not g3842 (n_1847, n2213);
  not g3843 (n_1848, n2219);
  and g3844 (n2221, n_1847, n_1848);
  not g3845 (n_1849, n2220);
  not g3846 (n_1850, n2221);
  and g3847 (n2222, n_1849, n_1850);
  and g3848 (n2223, n2190, n2222);
  not g3849 (n_1851, n2190);
  not g3850 (n_1852, n2222);
  and g3851 (n2224, n_1851, n_1852);
  not g3852 (n_1853, n2223);
  not g3853 (n_1854, n2224);
  and g3854 (n2225, n_1853, n_1854);
  and g3855 (n2226, n_1677, n_1703);
  and g3856 (n2227, \a[26] , \a[27] );
  and g3857 (n2228, n209, n2227);
  and g3858 (n2229, \a[8] , \a[27] );
  and g3859 (n2230, n1580, n2229);
  not g3860 (n_1855, n2228);
  not g3861 (n_1856, n2230);
  and g3862 (n2231, n_1855, n_1856);
  and g3863 (n2232, \a[4] , \a[26] );
  and g3864 (n2233, \a[8] , \a[22] );
  and g3865 (n2234, n2232, n2233);
  not g3866 (n_1857, n2231);
  not g3867 (n_1858, n2234);
  and g3868 (n2235, n_1857, n_1858);
  not g3869 (n_1859, n2235);
  and g3870 (n2236, n_1858, n_1859);
  not g3871 (n_1860, n2232);
  not g3872 (n_1861, n2233);
  and g3873 (n2237, n_1860, n_1861);
  not g3874 (n_1862, n2237);
  and g3875 (n2238, n2236, n_1862);
  and g3876 (n2239, \a[27] , n_1859);
  and g3877 (n2240, \a[3] , n2239);
  not g3878 (n_1863, n2238);
  not g3879 (n_1864, n2240);
  and g3880 (n2241, n_1863, n_1864);
  and g3881 (n2242, n335, n1666);
  and g3882 (n2243, n268, n1547);
  and g3883 (n2244, n332, n1904);
  not g3884 (n_1865, n2243);
  not g3885 (n_1866, n2244);
  and g3886 (n2245, n_1865, n_1866);
  not g3887 (n_1867, n2242);
  not g3888 (n_1868, n2245);
  and g3889 (n2246, n_1867, n_1868);
  not g3890 (n_1869, n2246);
  and g3891 (n2247, \a[25] , n_1869);
  and g3892 (n2248, \a[5] , n2247);
  and g3893 (n2249, n_1867, n_1869);
  and g3894 (n2250, \a[6] , \a[24] );
  and g3895 (n2251, \a[7] , \a[23] );
  not g3896 (n_1870, n2250);
  not g3897 (n_1871, n2251);
  and g3898 (n2252, n_1870, n_1871);
  not g3899 (n_1872, n2252);
  and g3900 (n2253, n2249, n_1872);
  not g3901 (n_1873, n2248);
  not g3902 (n_1874, n2253);
  and g3903 (n2254, n_1873, n_1874);
  not g3904 (n_1875, n2241);
  not g3905 (n_1876, n2254);
  and g3906 (n2255, n_1875, n_1876);
  not g3907 (n_1877, n2255);
  and g3908 (n2256, n_1875, n_1877);
  and g3909 (n2257, n_1876, n_1877);
  not g3910 (n_1878, n2256);
  not g3911 (n_1879, n2257);
  and g3912 (n2258, n_1878, n_1879);
  and g3913 (n2259, n602, n1149);
  and g3914 (n2260, n480, n1331);
  and g3915 (n2261, n723, n1490);
  not g3916 (n_1880, n2260);
  not g3917 (n_1881, n2261);
  and g3918 (n2262, n_1880, n_1881);
  not g3919 (n_1882, n2259);
  not g3920 (n_1883, n2262);
  and g3921 (n2263, n_1882, n_1883);
  not g3922 (n_1884, n2263);
  and g3923 (n2264, \a[20] , n_1884);
  and g3924 (n2265, \a[10] , n2264);
  and g3925 (n2266, \a[11] , \a[19] );
  and g3926 (n2267, \a[12] , \a[18] );
  not g3927 (n_1885, n2266);
  not g3928 (n_1886, n2267);
  and g3929 (n2268, n_1885, n_1886);
  and g3930 (n2269, n_1882, n_1884);
  not g3931 (n_1887, n2268);
  and g3932 (n2270, n_1887, n2269);
  not g3933 (n_1888, n2265);
  not g3934 (n_1889, n2270);
  and g3935 (n2271, n_1888, n_1889);
  not g3936 (n_1890, n2258);
  not g3937 (n_1891, n2271);
  and g3938 (n2272, n_1890, n_1891);
  not g3939 (n_1892, n2272);
  and g3940 (n2273, n_1890, n_1892);
  and g3941 (n2274, n_1891, n_1892);
  not g3942 (n_1893, n2273);
  not g3943 (n_1894, n2274);
  and g3944 (n2275, n_1893, n_1894);
  and g3945 (n2276, n_1715, n_1721);
  and g3946 (n2277, n2275, n2276);
  not g3947 (n_1895, n2275);
  not g3948 (n_1896, n2276);
  and g3949 (n2278, n_1895, n_1896);
  not g3950 (n_1897, n2277);
  not g3951 (n_1898, n2278);
  and g3952 (n2279, n_1897, n_1898);
  and g3953 (n2280, n_1682, n_1702);
  not g3954 (n_1899, n2280);
  and g3955 (n2281, n2279, n_1899);
  not g3956 (n_1900, n2279);
  and g3957 (n2282, n_1900, n2280);
  not g3958 (n_1901, n2281);
  not g3959 (n_1902, n2282);
  and g3960 (n2283, n_1901, n_1902);
  not g3961 (n_1903, n2226);
  and g3962 (n2284, n_1903, n2283);
  not g3963 (n_1904, n2283);
  and g3964 (n2285, n2226, n_1904);
  not g3965 (n_1905, n2284);
  not g3966 (n_1906, n2285);
  and g3967 (n2286, n_1905, n_1906);
  and g3968 (n2287, n2225, n2286);
  not g3969 (n_1907, n2225);
  not g3970 (n_1908, n2286);
  and g3971 (n2288, n_1907, n_1908);
  not g3972 (n_1909, n2287);
  not g3973 (n_1910, n2288);
  and g3974 (n2289, n_1909, n_1910);
  not g3975 (n_1911, n2164);
  and g3976 (n2290, n_1911, n2289);
  not g3977 (n_1912, n2289);
  and g3978 (n2291, n2164, n_1912);
  not g3979 (n_1913, n2290);
  not g3980 (n_1914, n2291);
  and g3981 (n2292, n_1913, n_1914);
  and g3982 (n2293, n_1790, n_1793);
  not g3983 (n_1915, n2293);
  and g3984 (n2294, n_1789, n_1915);
  not g3985 (n_1916, n2292);
  and g3986 (n2295, n_1916, n2294);
  not g3987 (n_1917, n2294);
  and g3988 (n2296, n2292, n_1917);
  not g3989 (n_1918, n2295);
  not g3990 (n_1919, n2296);
  and g3991 (\asquared[31] , n_1918, n_1919);
  and g3992 (n2298, n_1905, n_1909);
  and g3993 (n2299, n_1819, n_1853);
  and g3994 (n2300, n_1838, n_1849);
  and g3995 (n2301, \a[24] , \a[26] );
  and g3996 (n2302, n268, n2301);
  and g3997 (n2303, \a[23] , \a[26] );
  and g3998 (n2304, n354, n2303);
  and g3999 (n2305, n380, n1666);
  not g4000 (n_1920, n2304);
  not g4001 (n_1921, n2305);
  and g4002 (n2306, n_1920, n_1921);
  not g4003 (n_1922, n2302);
  not g4004 (n_1923, n2306);
  and g4005 (n2307, n_1922, n_1923);
  not g4006 (n_1924, n2307);
  and g4007 (n2308, n_1922, n_1924);
  and g4008 (n2309, \a[5] , \a[26] );
  and g4009 (n2310, \a[7] , \a[24] );
  not g4010 (n_1925, n2309);
  not g4011 (n_1926, n2310);
  and g4012 (n2311, n_1925, n_1926);
  not g4013 (n_1927, n2311);
  and g4014 (n2312, n2308, n_1927);
  and g4015 (n2313, \a[23] , n_1924);
  and g4016 (n2314, \a[8] , n2313);
  not g4017 (n_1928, n2312);
  not g4018 (n_1929, n2314);
  and g4019 (n2315, n_1928, n_1929);
  and g4020 (n2316, \a[14] , \a[17] );
  not g4021 (n_1930, n891);
  not g4022 (n_1931, n2316);
  and g4023 (n2317, n_1930, n_1931);
  and g4024 (n2318, n895, n1048);
  not g4025 (n_1932, n2318);
  not g4028 (n_1933, n2317);
  not g4030 (n_1934, n2321);
  and g4031 (n2322, \a[25] , n_1934);
  and g4032 (n2323, \a[6] , n2322);
  and g4033 (n2324, n_1932, n_1934);
  and g4034 (n2325, n_1933, n2324);
  not g4035 (n_1935, n2323);
  not g4036 (n_1936, n2325);
  and g4037 (n2326, n_1935, n_1936);
  not g4038 (n_1937, n2315);
  not g4039 (n_1938, n2326);
  and g4040 (n2327, n_1937, n_1938);
  not g4041 (n_1939, n2327);
  and g4042 (n2328, n_1937, n_1939);
  and g4043 (n2329, n_1938, n_1939);
  not g4044 (n_1940, n2328);
  not g4045 (n_1941, n2329);
  and g4046 (n2330, n_1940, n_1941);
  and g4047 (n2331, \a[27] , \a[28] );
  and g4048 (n2332, n209, n2331);
  and g4049 (n2333, n252, n2041);
  and g4050 (n2334, \a[28] , \a[29] );
  and g4051 (n2335, n218, n2334);
  not g4052 (n_1942, n2333);
  not g4053 (n_1943, n2335);
  and g4054 (n2336, n_1942, n_1943);
  not g4055 (n_1944, n2332);
  not g4056 (n_1945, n2336);
  and g4057 (n2337, n_1944, n_1945);
  not g4058 (n_1946, n2337);
  and g4059 (n2338, \a[29] , n_1946);
  and g4060 (n2339, \a[2] , n2338);
  and g4061 (n2340, \a[3] , \a[28] );
  and g4062 (n2341, \a[4] , \a[27] );
  not g4063 (n_1947, n2340);
  not g4064 (n_1948, n2341);
  and g4065 (n2342, n_1947, n_1948);
  and g4066 (n2343, n_1944, n_1946);
  not g4067 (n_1949, n2342);
  and g4068 (n2344, n_1949, n2343);
  not g4069 (n_1950, n2339);
  not g4070 (n_1951, n2344);
  and g4071 (n2345, n_1950, n_1951);
  not g4072 (n_1952, n2330);
  not g4073 (n_1953, n2345);
  and g4074 (n2346, n_1952, n_1953);
  not g4075 (n_1954, n2346);
  and g4076 (n2347, n_1952, n_1954);
  and g4077 (n2348, n_1953, n_1954);
  not g4078 (n_1955, n2347);
  not g4079 (n_1956, n2348);
  and g4080 (n2349, n_1955, n_1956);
  and g4081 (n2350, \a[22] , \a[31] );
  and g4082 (n2351, n350, n2350);
  and g4083 (n2352, \a[10] , \a[31] );
  and g4084 (n2353, n1199, n2352);
  and g4085 (n2354, n484, n1574);
  not g4086 (n_1958, n2353);
  not g4087 (n_1959, n2354);
  and g4088 (n2355, n_1958, n_1959);
  not g4089 (n_1960, n2351);
  not g4090 (n_1961, n2355);
  and g4091 (n2356, n_1960, n_1961);
  not g4092 (n_1962, n2356);
  and g4093 (n2357, n_1960, n_1962);
  and g4094 (n2358, \a[0] , \a[31] );
  and g4095 (n2359, \a[9] , \a[22] );
  not g4096 (n_1963, n2358);
  not g4097 (n_1964, n2359);
  and g4098 (n2360, n_1963, n_1964);
  not g4099 (n_1965, n2360);
  and g4100 (n2361, n2357, n_1965);
  and g4101 (n2362, \a[21] , n_1962);
  and g4102 (n2363, \a[10] , n2362);
  not g4103 (n_1966, n2361);
  not g4104 (n_1967, n2363);
  and g4105 (n2364, n_1966, n_1967);
  and g4106 (n2365, n_1797, n_1805);
  and g4107 (n2366, n748, n1149);
  and g4108 (n2367, n818, n1331);
  and g4109 (n2368, n602, n1490);
  not g4110 (n_1968, n2367);
  not g4111 (n_1969, n2368);
  and g4112 (n2369, n_1968, n_1969);
  not g4113 (n_1970, n2366);
  not g4114 (n_1971, n2369);
  and g4115 (n2370, n_1970, n_1971);
  not g4116 (n_1972, n2370);
  and g4117 (n2371, \a[20] , n_1972);
  and g4118 (n2372, \a[11] , n2371);
  and g4119 (n2373, n_1970, n_1972);
  and g4120 (n2374, \a[12] , \a[19] );
  and g4121 (n2375, \a[13] , \a[18] );
  not g4122 (n_1973, n2374);
  not g4123 (n_1974, n2375);
  and g4124 (n2376, n_1973, n_1974);
  not g4125 (n_1975, n2376);
  and g4126 (n2377, n2373, n_1975);
  not g4127 (n_1976, n2372);
  not g4128 (n_1977, n2377);
  and g4129 (n2378, n_1976, n_1977);
  not g4130 (n_1978, n2365);
  not g4131 (n_1979, n2378);
  and g4132 (n2379, n_1978, n_1979);
  not g4133 (n_1980, n2379);
  and g4134 (n2380, n_1978, n_1980);
  and g4135 (n2381, n_1979, n_1980);
  not g4136 (n_1981, n2380);
  not g4137 (n_1982, n2381);
  and g4138 (n2382, n_1981, n_1982);
  not g4139 (n_1983, n2364);
  not g4140 (n_1984, n2382);
  and g4141 (n2383, n_1983, n_1984);
  and g4142 (n2384, n2364, n_1982);
  and g4143 (n2385, n_1981, n2384);
  not g4144 (n_1985, n2383);
  not g4145 (n_1986, n2385);
  and g4146 (n2386, n_1985, n_1986);
  not g4147 (n_1987, n2349);
  and g4148 (n2387, n_1987, n2386);
  not g4149 (n_1988, n2386);
  and g4150 (n2388, n2349, n_1988);
  not g4151 (n_1989, n2387);
  not g4152 (n_1990, n2388);
  and g4153 (n2389, n_1989, n_1990);
  not g4154 (n_1991, n2300);
  and g4155 (n2390, n_1991, n2389);
  not g4156 (n_1992, n2389);
  and g4157 (n2391, n2300, n_1992);
  not g4158 (n_1993, n2390);
  not g4159 (n_1994, n2391);
  and g4160 (n2392, n_1993, n_1994);
  not g4161 (n_1995, n2299);
  and g4162 (n2393, n_1995, n2392);
  not g4163 (n_1996, n2392);
  and g4164 (n2394, n2299, n_1996);
  not g4165 (n_1997, n2393);
  not g4166 (n_1998, n2394);
  and g4167 (n2395, n_1997, n_1998);
  and g4168 (n2396, n_1898, n_1901);
  and g4169 (n2397, n_1823, n_1832);
  and g4170 (n2398, n_1842, n_1846);
  and g4171 (n2399, n2397, n2398);
  not g4172 (n_1999, n2397);
  not g4173 (n_2000, n2398);
  and g4174 (n2400, n_1999, n_2000);
  not g4175 (n_2001, n2399);
  not g4176 (n_2002, n2400);
  and g4177 (n2401, n_2001, n_2002);
  and g4178 (n2402, \a[1] , \a[30] );
  and g4179 (n2403, \a[16] , n2402);
  not g4180 (n_2003, \a[16] );
  not g4181 (n_2004, n2402);
  and g4182 (n2404, n_2003, n_2004);
  not g4183 (n_2005, n2403);
  not g4184 (n_2006, n2404);
  and g4185 (n2405, n_2005, n_2006);
  and g4186 (n2406, n2171, n2405);
  not g4187 (n_2007, n2405);
  and g4188 (n2407, n_1800, n_2007);
  not g4189 (n_2008, n2406);
  not g4190 (n_2009, n2407);
  and g4191 (n2408, n_2008, n_2009);
  not g4192 (n_2010, n2249);
  and g4193 (n2409, n_2010, n2408);
  not g4194 (n_2011, n2408);
  and g4195 (n2410, n2249, n_2011);
  not g4196 (n_2012, n2409);
  not g4197 (n_2013, n2410);
  and g4198 (n2411, n_2012, n_2013);
  and g4199 (n2412, n2401, n2411);
  not g4200 (n_2014, n2401);
  not g4201 (n_2015, n2411);
  and g4202 (n2413, n_2014, n_2015);
  not g4203 (n_2016, n2412);
  not g4204 (n_2017, n2413);
  and g4205 (n2414, n_2016, n_2017);
  not g4206 (n_2018, n2414);
  and g4207 (n2415, n2396, n_2018);
  not g4208 (n_2019, n2396);
  and g4209 (n2416, n_2019, n2414);
  not g4210 (n_2020, n2415);
  not g4211 (n_2021, n2416);
  and g4212 (n2417, n_2020, n_2021);
  and g4213 (n2418, n2203, n2236);
  not g4214 (n_2022, n2203);
  not g4215 (n_2023, n2236);
  and g4216 (n2419, n_2022, n_2023);
  not g4217 (n_2024, n2418);
  not g4218 (n_2025, n2419);
  and g4219 (n2420, n_2024, n_2025);
  not g4220 (n_2026, n2420);
  and g4221 (n2421, n2269, n_2026);
  not g4222 (n_2027, n2269);
  and g4223 (n2422, n_2027, n2420);
  not g4224 (n_2028, n2421);
  not g4225 (n_2029, n2422);
  and g4226 (n2423, n_2028, n_2029);
  and g4227 (n2424, n_1877, n_1892);
  not g4228 (n_2030, n2423);
  and g4229 (n2425, n_2030, n2424);
  not g4230 (n_2031, n2424);
  and g4231 (n2426, n2423, n_2031);
  not g4232 (n_2032, n2425);
  not g4233 (n_2033, n2426);
  and g4234 (n2427, n_2032, n_2033);
  and g4235 (n2428, n_1811, n_1815);
  not g4236 (n_2034, n2427);
  and g4237 (n2429, n_2034, n2428);
  not g4238 (n_2035, n2428);
  and g4239 (n2430, n2427, n_2035);
  not g4240 (n_2036, n2429);
  not g4241 (n_2037, n2430);
  and g4242 (n2431, n_2036, n_2037);
  and g4243 (n2432, n2417, n2431);
  not g4244 (n_2038, n2417);
  not g4245 (n_2039, n2431);
  and g4246 (n2433, n_2038, n_2039);
  not g4247 (n_2040, n2432);
  not g4248 (n_2041, n2433);
  and g4249 (n2434, n_2040, n_2041);
  and g4250 (n2435, n2395, n2434);
  not g4251 (n_2042, n2395);
  not g4252 (n_2043, n2434);
  and g4253 (n2436, n_2042, n_2043);
  not g4254 (n_2044, n2435);
  not g4255 (n_2045, n2436);
  and g4256 (n2437, n_2044, n_2045);
  not g4257 (n_2046, n2298);
  and g4258 (n2438, n_2046, n2437);
  not g4259 (n_2047, n2437);
  and g4260 (n2439, n2298, n_2047);
  not g4261 (n_2048, n2438);
  not g4262 (n_2049, n2439);
  and g4263 (n2440, n_2048, n_2049);
  and g4264 (n2441, n_1914, n_1917);
  not g4265 (n_2050, n2441);
  and g4266 (n2442, n_1913, n_2050);
  not g4267 (n_2051, n2440);
  and g4268 (n2443, n_2051, n2442);
  not g4269 (n_2052, n2442);
  and g4270 (n2444, n2440, n_2052);
  not g4271 (n_2053, n2443);
  not g4272 (n_2054, n2444);
  and g4273 (\asquared[32] , n_2053, n_2054);
  and g4274 (n2446, n_2049, n_2052);
  not g4275 (n_2055, n2446);
  and g4276 (n2447, n_2048, n_2055);
  and g4277 (n2448, n_1997, n_2044);
  and g4278 (n2449, n_2021, n_2040);
  and g4279 (n2450, n_2033, n_2037);
  and g4280 (n2451, \a[5] , \a[27] );
  and g4281 (n2452, \a[4] , \a[28] );
  not g4282 (n_2056, n2451);
  not g4283 (n_2057, n2452);
  and g4284 (n2453, n_2056, n_2057);
  and g4285 (n2454, n226, n2331);
  not g4286 (n_2058, n2454);
  not g4289 (n_2059, n2453);
  not g4291 (n_2060, n2457);
  and g4292 (n2458, n_2058, n_2060);
  and g4293 (n2459, n_2059, n2458);
  and g4294 (n2460, \a[23] , n_2060);
  and g4295 (n2461, \a[9] , n2460);
  not g4296 (n_2061, n2459);
  not g4297 (n_2062, n2461);
  and g4298 (n2462, n_2061, n_2062);
  and g4299 (n2463, \a[25] , \a[26] );
  and g4300 (n2464, n335, n2463);
  and g4301 (n2465, n312, n2301);
  and g4302 (n2466, n380, n1904);
  not g4303 (n_2063, n2465);
  not g4304 (n_2064, n2466);
  and g4305 (n2467, n_2063, n_2064);
  not g4306 (n_2065, n2464);
  not g4307 (n_2066, n2467);
  and g4308 (n2468, n_2065, n_2066);
  not g4309 (n_2067, n2468);
  and g4310 (n2469, \a[24] , n_2067);
  and g4311 (n2470, \a[8] , n2469);
  and g4312 (n2471, n_2065, n_2067);
  and g4313 (n2472, \a[6] , \a[26] );
  and g4314 (n2473, \a[7] , \a[25] );
  not g4315 (n_2068, n2472);
  not g4316 (n_2069, n2473);
  and g4317 (n2474, n_2068, n_2069);
  not g4318 (n_2070, n2474);
  and g4319 (n2475, n2471, n_2070);
  not g4320 (n_2071, n2470);
  not g4321 (n_2072, n2475);
  and g4322 (n2476, n_2071, n_2072);
  not g4323 (n_2073, n2462);
  not g4324 (n_2074, n2476);
  and g4325 (n2477, n_2073, n_2074);
  not g4326 (n_2075, n2477);
  and g4327 (n2478, n_2073, n_2075);
  and g4328 (n2479, n_2074, n_2075);
  not g4329 (n_2076, n2478);
  not g4330 (n_2077, n2479);
  and g4331 (n2480, n_2076, n_2077);
  and g4332 (n2481, n_2008, n_2012);
  and g4333 (n2482, n2480, n2481);
  not g4334 (n_2078, n2480);
  not g4335 (n_2079, n2481);
  and g4336 (n2483, n_2078, n_2079);
  not g4337 (n_2080, n2482);
  not g4338 (n_2081, n2483);
  and g4339 (n2484, n_2080, n_2081);
  and g4340 (n2485, \a[0] , \a[32] );
  and g4341 (n2486, \a[2] , \a[30] );
  not g4342 (n_2083, n2485);
  not g4343 (n_2084, n2486);
  and g4344 (n2487, n_2083, n_2084);
  and g4345 (n2488, \a[30] , \a[32] );
  and g4346 (n2489, n196, n2488);
  not g4347 (n_2085, n2487);
  not g4348 (n_2086, n2489);
  and g4349 (n2490, n_2085, n_2086);
  and g4350 (n2491, n2403, n2490);
  not g4351 (n_2087, n2491);
  and g4352 (n2492, n_2086, n_2087);
  and g4353 (n2493, n_2085, n2492);
  and g4354 (n2494, n2403, n_2087);
  not g4355 (n_2088, n2493);
  not g4356 (n_2089, n2494);
  and g4357 (n2495, n_2088, n_2089);
  and g4358 (n2496, n748, n1490);
  and g4359 (n2497, n818, n1492);
  and g4360 (n2498, n602, n1494);
  not g4361 (n_2090, n2497);
  not g4362 (n_2091, n2498);
  and g4363 (n2499, n_2090, n_2091);
  not g4364 (n_2092, n2496);
  not g4365 (n_2093, n2499);
  and g4366 (n2500, n_2092, n_2093);
  not g4367 (n_2094, n2500);
  and g4368 (n2501, \a[21] , n_2094);
  and g4369 (n2502, \a[11] , n2501);
  and g4370 (n2503, n_2092, n_2094);
  and g4371 (n2504, \a[12] , \a[20] );
  and g4372 (n2505, \a[13] , \a[19] );
  not g4373 (n_2095, n2504);
  not g4374 (n_2096, n2505);
  and g4375 (n2506, n_2095, n_2096);
  not g4376 (n_2097, n2506);
  and g4377 (n2507, n2503, n_2097);
  not g4378 (n_2098, n2502);
  not g4379 (n_2099, n2507);
  and g4380 (n2508, n_2098, n_2099);
  not g4381 (n_2100, n2495);
  not g4382 (n_2101, n2508);
  and g4383 (n2509, n_2100, n_2101);
  not g4384 (n_2102, n2509);
  and g4385 (n2510, n_2100, n_2102);
  and g4386 (n2511, n_2101, n_2102);
  not g4387 (n_2103, n2510);
  not g4388 (n_2104, n2511);
  and g4389 (n2512, n_2103, n_2104);
  and g4390 (n2513, \a[3] , \a[29] );
  and g4391 (n2514, \a[10] , \a[22] );
  not g4392 (n_2105, n2513);
  not g4393 (n_2106, n2514);
  and g4394 (n2515, n_2105, n_2106);
  and g4395 (n2516, n2513, n2514);
  not g4396 (n_2107, n2516);
  not g4399 (n_2108, n2515);
  not g4401 (n_2109, n2519);
  and g4402 (n2520, \a[18] , n_2109);
  and g4403 (n2521, \a[14] , n2520);
  and g4404 (n2522, n_2107, n_2109);
  and g4405 (n2523, n_2108, n2522);
  not g4406 (n_2110, n2521);
  not g4407 (n_2111, n2523);
  and g4408 (n2524, n_2110, n_2111);
  not g4409 (n_2112, n2512);
  not g4410 (n_2113, n2524);
  and g4411 (n2525, n_2112, n_2113);
  not g4412 (n_2114, n2525);
  and g4413 (n2526, n_2112, n_2114);
  and g4414 (n2527, n_2113, n_2114);
  not g4415 (n_2115, n2526);
  not g4416 (n_2116, n2527);
  and g4417 (n2528, n_2115, n_2116);
  not g4418 (n_2117, n2484);
  and g4419 (n2529, n_2117, n2528);
  not g4420 (n_2118, n2528);
  and g4421 (n2530, n2484, n_2118);
  not g4422 (n_2119, n2529);
  not g4423 (n_2120, n2530);
  and g4424 (n2531, n_2119, n_2120);
  not g4425 (n_2121, n2450);
  and g4426 (n2532, n_2121, n2531);
  not g4427 (n_2122, n2531);
  and g4428 (n2533, n2450, n_2122);
  not g4429 (n_2123, n2532);
  not g4430 (n_2124, n2533);
  and g4431 (n2534, n_2123, n_2124);
  not g4432 (n_2125, n2449);
  and g4433 (n2535, n_2125, n2534);
  not g4434 (n_2126, n2534);
  and g4435 (n2536, n2449, n_2126);
  not g4436 (n_2127, n2535);
  not g4437 (n_2128, n2536);
  and g4438 (n2537, n_2127, n_2128);
  and g4439 (n2538, n_2002, n_2016);
  and g4440 (n2539, n2357, n2373);
  not g4441 (n_2129, n2357);
  not g4442 (n_2130, n2373);
  and g4443 (n2540, n_2129, n_2130);
  not g4444 (n_2131, n2539);
  not g4445 (n_2132, n2540);
  and g4446 (n2541, n_2131, n_2132);
  not g4447 (n_2133, n2541);
  and g4448 (n2542, n2343, n_2133);
  not g4449 (n_2134, n2343);
  and g4450 (n2543, n_2134, n2541);
  not g4451 (n_2135, n2542);
  not g4452 (n_2136, n2543);
  and g4453 (n2544, n_2135, n_2136);
  and g4454 (n2545, \a[1] , \a[31] );
  not g4455 (n_2137, n993);
  not g4456 (n_2138, n2545);
  and g4457 (n2546, n_2137, n_2138);
  and g4458 (n2547, n993, n2545);
  not g4459 (n_2139, n2546);
  not g4460 (n_2140, n2547);
  and g4461 (n2548, n_2139, n_2140);
  not g4462 (n_2141, n2548);
  and g4463 (n2549, n2324, n_2141);
  not g4464 (n_2142, n2324);
  and g4465 (n2550, n_2142, n2548);
  not g4466 (n_2143, n2549);
  not g4467 (n_2144, n2550);
  and g4468 (n2551, n_2143, n_2144);
  not g4469 (n_2145, n2308);
  and g4470 (n2552, n_2145, n2551);
  not g4471 (n_2146, n2551);
  and g4472 (n2553, n2308, n_2146);
  not g4473 (n_2147, n2552);
  not g4474 (n_2148, n2553);
  and g4475 (n2554, n_2147, n_2148);
  and g4476 (n2555, n2544, n2554);
  not g4477 (n_2149, n2544);
  not g4478 (n_2150, n2554);
  and g4479 (n2556, n_2149, n_2150);
  not g4480 (n_2151, n2555);
  not g4481 (n_2152, n2556);
  and g4482 (n2557, n_2151, n_2152);
  not g4483 (n_2153, n2557);
  and g4484 (n2558, n2538, n_2153);
  not g4485 (n_2154, n2538);
  and g4486 (n2559, n_2154, n2557);
  not g4487 (n_2155, n2558);
  not g4488 (n_2156, n2559);
  and g4489 (n2560, n_2155, n_2156);
  and g4490 (n2561, n_1980, n_1985);
  and g4491 (n2562, n_2025, n_2029);
  and g4492 (n2563, n2561, n2562);
  not g4493 (n_2157, n2561);
  not g4494 (n_2158, n2562);
  and g4495 (n2564, n_2157, n_2158);
  not g4496 (n_2159, n2563);
  not g4497 (n_2160, n2564);
  and g4498 (n2565, n_2159, n_2160);
  and g4499 (n2566, n_1939, n_1954);
  not g4500 (n_2161, n2565);
  and g4501 (n2567, n_2161, n2566);
  not g4502 (n_2162, n2566);
  and g4503 (n2568, n2565, n_2162);
  not g4504 (n_2163, n2567);
  not g4505 (n_2164, n2568);
  and g4506 (n2569, n_2163, n_2164);
  and g4507 (n2570, n_1989, n_1993);
  not g4508 (n_2165, n2569);
  and g4509 (n2571, n_2165, n2570);
  not g4510 (n_2166, n2570);
  and g4511 (n2572, n2569, n_2166);
  not g4512 (n_2167, n2571);
  not g4513 (n_2168, n2572);
  and g4514 (n2573, n_2167, n_2168);
  and g4515 (n2574, n2560, n2573);
  not g4516 (n_2169, n2560);
  not g4517 (n_2170, n2573);
  and g4518 (n2575, n_2169, n_2170);
  not g4519 (n_2171, n2574);
  not g4520 (n_2172, n2575);
  and g4521 (n2576, n_2171, n_2172);
  and g4522 (n2577, n2537, n2576);
  not g4523 (n_2173, n2537);
  not g4524 (n_2174, n2576);
  and g4525 (n2578, n_2173, n_2174);
  not g4526 (n_2175, n2577);
  not g4527 (n_2176, n2578);
  and g4528 (n2579, n_2175, n_2176);
  not g4529 (n_2177, n2448);
  and g4530 (n2580, n_2177, n2579);
  not g4531 (n_2178, n2579);
  and g4532 (n2581, n2448, n_2178);
  not g4533 (n_2179, n2580);
  not g4534 (n_2180, n2581);
  and g4535 (n2582, n_2179, n_2180);
  not g4536 (n_2181, n2447);
  and g4537 (n2583, n_2181, n2582);
  not g4538 (n_2182, n2582);
  and g4539 (n2584, n2447, n_2182);
  not g4540 (n_2183, n2583);
  not g4541 (n_2184, n2584);
  and g4542 (\asquared[33] , n_2183, n_2184);
  and g4543 (n2586, n2492, n2503);
  not g4544 (n_2185, n2492);
  not g4545 (n_2186, n2503);
  and g4546 (n2587, n_2185, n_2186);
  not g4547 (n_2187, n2586);
  not g4548 (n_2188, n2587);
  and g4549 (n2588, n_2187, n_2188);
  not g4550 (n_2189, n2588);
  and g4551 (n2589, n2522, n_2189);
  not g4552 (n_2190, n2522);
  and g4553 (n2590, n_2190, n2588);
  not g4554 (n_2191, n2589);
  not g4555 (n_2192, n2590);
  and g4556 (n2591, n_2191, n_2192);
  and g4557 (n2592, n2458, n2471);
  not g4558 (n_2193, n2458);
  not g4559 (n_2194, n2471);
  and g4560 (n2593, n_2193, n_2194);
  not g4561 (n_2195, n2592);
  not g4562 (n_2196, n2593);
  and g4563 (n2594, n_2195, n_2196);
  and g4564 (n2595, \a[22] , \a[33] );
  and g4565 (n2596, n449, n2595);
  and g4566 (n2597, n544, n2350);
  and g4567 (n2598, \a[31] , \a[33] );
  and g4568 (n2599, n196, n2598);
  not g4569 (n_2198, n2597);
  not g4570 (n_2199, n2599);
  and g4571 (n2600, n_2198, n_2199);
  not g4572 (n_2200, n2596);
  not g4573 (n_2201, n2600);
  and g4574 (n2601, n_2200, n_2201);
  not g4575 (n_2202, n2601);
  and g4576 (n2602, \a[31] , n_2202);
  and g4577 (n2603, \a[2] , n2602);
  and g4578 (n2604, n_2200, n_2202);
  and g4579 (n2605, \a[0] , \a[33] );
  and g4580 (n2606, \a[11] , \a[22] );
  not g4581 (n_2203, n2605);
  not g4582 (n_2204, n2606);
  and g4583 (n2607, n_2203, n_2204);
  not g4584 (n_2205, n2607);
  and g4585 (n2608, n2604, n_2205);
  not g4586 (n_2206, n2603);
  not g4587 (n_2207, n2608);
  and g4588 (n2609, n_2206, n_2207);
  not g4589 (n_2208, n2609);
  and g4590 (n2610, n2594, n_2208);
  not g4591 (n_2209, n2610);
  and g4592 (n2611, n2594, n_2209);
  and g4593 (n2612, n_2208, n_2209);
  not g4594 (n_2210, n2611);
  not g4595 (n_2211, n2612);
  and g4596 (n2613, n_2210, n_2211);
  not g4597 (n_2212, n2591);
  and g4598 (n2614, n_2212, n2613);
  not g4599 (n_2213, n2613);
  and g4600 (n2615, n2591, n_2213);
  not g4601 (n_2214, n2614);
  not g4602 (n_2215, n2615);
  and g4603 (n2616, n_2214, n_2215);
  and g4604 (n2617, \a[29] , \a[30] );
  and g4605 (n2618, n209, n2617);
  and g4606 (n2619, \a[24] , \a[30] );
  and g4607 (n2620, n479, n2619);
  not g4608 (n_2216, n2618);
  not g4609 (n_2217, n2620);
  and g4610 (n2621, n_2216, n_2217);
  and g4611 (n2622, \a[4] , \a[29] );
  and g4612 (n2623, \a[9] , \a[24] );
  and g4613 (n2624, n2622, n2623);
  not g4614 (n_2218, n2621);
  not g4615 (n_2219, n2624);
  and g4616 (n2625, n_2218, n_2219);
  not g4617 (n_2220, n2625);
  and g4618 (n2626, n_2219, n_2220);
  not g4619 (n_2221, n2622);
  not g4620 (n_2222, n2623);
  and g4621 (n2627, n_2221, n_2222);
  not g4622 (n_2223, n2627);
  and g4623 (n2628, n2626, n_2223);
  and g4624 (n2629, \a[30] , n_2220);
  and g4625 (n2630, \a[3] , n2629);
  not g4626 (n_2224, n2628);
  not g4627 (n_2225, n2630);
  and g4628 (n2631, n_2224, n_2225);
  and g4629 (n2632, \a[5] , \a[28] );
  and g4630 (n2633, \a[25] , \a[27] );
  and g4631 (n2634, n312, n2633);
  and g4632 (n2635, n332, n2331);
  and g4633 (n2636, \a[8] , \a[25] );
  and g4634 (n2637, n2632, n2636);
  not g4635 (n_2226, n2635);
  not g4636 (n_2227, n2637);
  and g4637 (n2638, n_2226, n_2227);
  not g4638 (n_2228, n2634);
  not g4639 (n_2229, n2638);
  and g4640 (n2639, n_2228, n_2229);
  not g4641 (n_2230, n2639);
  and g4642 (n2640, n2632, n_2230);
  and g4643 (n2641, \a[6] , \a[27] );
  not g4644 (n_2231, n2636);
  not g4645 (n_2232, n2641);
  and g4646 (n2642, n_2231, n_2232);
  and g4647 (n2643, n_2228, n_2230);
  not g4648 (n_2233, n2642);
  and g4649 (n2644, n_2233, n2643);
  not g4650 (n_2234, n2640);
  not g4651 (n_2235, n2644);
  and g4652 (n2645, n_2234, n_2235);
  not g4653 (n_2236, n2631);
  not g4654 (n_2237, n2645);
  and g4655 (n2646, n_2236, n_2237);
  not g4656 (n_2238, n2646);
  and g4657 (n2647, n_2236, n_2238);
  and g4658 (n2648, n_2237, n_2238);
  not g4659 (n_2239, n2647);
  not g4660 (n_2240, n2648);
  and g4661 (n2649, n_2239, n_2240);
  and g4662 (n2650, \a[15] , \a[18] );
  not g4663 (n_2241, n1048);
  not g4664 (n_2242, n2650);
  and g4665 (n2651, n_2241, n_2242);
  and g4666 (n2652, n891, n1052);
  not g4667 (n_2243, n2652);
  not g4670 (n_2244, n2651);
  not g4672 (n_2245, n2655);
  and g4673 (n2656, \a[26] , n_2245);
  and g4674 (n2657, \a[7] , n2656);
  and g4675 (n2658, n_2243, n_2245);
  and g4676 (n2659, n_2244, n2658);
  not g4677 (n_2246, n2657);
  not g4678 (n_2247, n2659);
  and g4679 (n2660, n_2246, n_2247);
  not g4680 (n_2248, n2649);
  not g4681 (n_2249, n2660);
  and g4682 (n2661, n_2248, n_2249);
  not g4683 (n_2250, n2661);
  and g4684 (n2662, n_2248, n_2250);
  and g4685 (n2663, n_2249, n_2250);
  not g4686 (n_2251, n2662);
  not g4687 (n_2252, n2663);
  and g4688 (n2664, n_2251, n_2252);
  and g4689 (n2665, n2616, n2664);
  not g4690 (n_2253, n2616);
  not g4691 (n_2254, n2664);
  and g4692 (n2666, n_2253, n_2254);
  not g4693 (n_2255, n2665);
  not g4694 (n_2256, n2666);
  and g4695 (n2667, n_2255, n_2256);
  and g4696 (n2668, n_2132, n_2136);
  and g4697 (n2669, n_2102, n_2114);
  and g4698 (n2670, n2668, n2669);
  not g4699 (n_2257, n2668);
  not g4700 (n_2258, n2669);
  and g4701 (n2671, n_2257, n_2258);
  not g4702 (n_2259, n2670);
  not g4703 (n_2260, n2671);
  and g4704 (n2672, n_2259, n_2260);
  and g4705 (n2673, n_2075, n_2081);
  not g4706 (n_2261, n2672);
  and g4707 (n2674, n_2261, n2673);
  not g4708 (n_2262, n2673);
  and g4709 (n2675, n2672, n_2262);
  not g4710 (n_2263, n2674);
  not g4711 (n_2264, n2675);
  and g4712 (n2676, n_2263, n_2264);
  and g4713 (n2677, n_2120, n_2123);
  not g4714 (n_2265, n2677);
  and g4715 (n2678, n2676, n_2265);
  not g4716 (n_2266, n2676);
  and g4717 (n2679, n_2266, n2677);
  not g4718 (n_2267, n2678);
  not g4719 (n_2268, n2679);
  and g4720 (n2680, n_2267, n_2268);
  not g4721 (n_2269, n2667);
  and g4722 (n2681, n_2269, n2680);
  not g4723 (n_2270, n2680);
  and g4724 (n2682, n2667, n_2270);
  not g4725 (n_2271, n2681);
  not g4726 (n_2272, n2682);
  and g4727 (n2683, n_2271, n_2272);
  and g4728 (n2684, \a[10] , \a[23] );
  not g4729 (n_2273, n2684);
  and g4730 (n2685, n_2140, n_2273);
  and g4731 (n2686, n2547, n2684);
  and g4732 (n2687, \a[1] , \a[32] );
  not g4733 (n_2274, n2687);
  and g4734 (n2688, \a[17] , n_2274);
  not g4735 (n_2275, \a[17] );
  and g4736 (n2689, n_2275, n2687);
  not g4737 (n_2276, n2688);
  not g4738 (n_2277, n2689);
  and g4739 (n2690, n_2276, n_2277);
  not g4740 (n_2278, n2686);
  not g4741 (n_2279, n2690);
  and g4742 (n2691, n_2278, n_2279);
  not g4743 (n_2280, n2685);
  and g4744 (n2692, n_2280, n2691);
  not g4745 (n_2281, n2692);
  and g4746 (n2693, n_2278, n_2281);
  and g4747 (n2694, n_2280, n2693);
  and g4748 (n2695, n_2279, n_2281);
  not g4749 (n_2282, n2694);
  not g4750 (n_2283, n2695);
  and g4751 (n2696, n_2282, n_2283);
  and g4752 (n2697, n745, n1490);
  and g4753 (n2698, n606, n1492);
  and g4754 (n2699, n748, n1494);
  not g4755 (n_2284, n2698);
  not g4756 (n_2285, n2699);
  and g4757 (n2700, n_2284, n_2285);
  not g4758 (n_2286, n2697);
  not g4759 (n_2287, n2700);
  and g4760 (n2701, n_2286, n_2287);
  not g4761 (n_2288, n2701);
  and g4762 (n2702, \a[21] , n_2288);
  and g4763 (n2703, \a[12] , n2702);
  and g4764 (n2704, n_2286, n_2288);
  and g4765 (n2705, \a[13] , \a[20] );
  and g4766 (n2706, \a[14] , \a[19] );
  not g4767 (n_2289, n2705);
  not g4768 (n_2290, n2706);
  and g4769 (n2707, n_2289, n_2290);
  not g4770 (n_2291, n2707);
  and g4771 (n2708, n2704, n_2291);
  not g4772 (n_2292, n2703);
  not g4773 (n_2293, n2708);
  and g4774 (n2709, n_2292, n_2293);
  not g4775 (n_2294, n2696);
  not g4776 (n_2295, n2709);
  and g4777 (n2710, n_2294, n_2295);
  not g4778 (n_2296, n2710);
  and g4779 (n2711, n_2294, n_2296);
  and g4780 (n2712, n_2295, n_2296);
  not g4781 (n_2297, n2711);
  not g4782 (n_2298, n2712);
  and g4783 (n2713, n_2297, n_2298);
  and g4784 (n2714, n_2144, n_2147);
  and g4785 (n2715, n2713, n2714);
  not g4786 (n_2299, n2713);
  not g4787 (n_2300, n2714);
  and g4788 (n2716, n_2299, n_2300);
  not g4789 (n_2301, n2715);
  not g4790 (n_2302, n2716);
  and g4791 (n2717, n_2301, n_2302);
  and g4792 (n2718, n_2160, n_2164);
  not g4793 (n_2303, n2717);
  and g4794 (n2719, n_2303, n2718);
  not g4795 (n_2304, n2718);
  and g4796 (n2720, n2717, n_2304);
  not g4797 (n_2305, n2719);
  not g4798 (n_2306, n2720);
  and g4799 (n2721, n_2305, n_2306);
  and g4800 (n2722, n_2151, n_2156);
  not g4801 (n_2307, n2721);
  and g4802 (n2723, n_2307, n2722);
  not g4803 (n_2308, n2722);
  and g4804 (n2724, n2721, n_2308);
  not g4805 (n_2309, n2723);
  not g4806 (n_2310, n2724);
  and g4807 (n2725, n_2309, n_2310);
  and g4808 (n2726, n_2168, n_2171);
  not g4809 (n_2311, n2726);
  and g4810 (n2727, n2725, n_2311);
  not g4811 (n_2312, n2725);
  and g4812 (n2728, n_2312, n2726);
  not g4813 (n_2313, n2727);
  not g4814 (n_2314, n2728);
  and g4815 (n2729, n_2313, n_2314);
  and g4816 (n2730, n2683, n2729);
  not g4817 (n_2315, n2683);
  not g4818 (n_2316, n2729);
  and g4819 (n2731, n_2315, n_2316);
  not g4820 (n_2317, n2730);
  not g4821 (n_2318, n2731);
  and g4822 (n2732, n_2317, n_2318);
  and g4823 (n2733, n_2127, n_2175);
  not g4824 (n_2319, n2732);
  and g4825 (n2734, n_2319, n2733);
  not g4826 (n_2320, n2733);
  and g4827 (n2735, n2732, n_2320);
  not g4828 (n_2321, n2734);
  not g4829 (n_2322, n2735);
  and g4830 (n2736, n_2321, n_2322);
  and g4831 (n2737, n_2181, n_2180);
  not g4832 (n_2323, n2737);
  and g4833 (n2738, n_2179, n_2323);
  not g4834 (n_2324, n2736);
  and g4835 (n2739, n_2324, n2738);
  not g4836 (n_2325, n2738);
  and g4837 (n2740, n2736, n_2325);
  not g4838 (n_2326, n2739);
  not g4839 (n_2327, n2740);
  and g4840 (\asquared[34] , n_2326, n_2327);
  and g4841 (n2742, n_2321, n_2325);
  not g4842 (n_2328, n2742);
  and g4843 (n2743, n_2322, n_2328);
  and g4844 (n2744, n_2313, n_2317);
  and g4845 (n2745, n2693, n2704);
  not g4846 (n_2329, n2693);
  not g4847 (n_2330, n2704);
  and g4848 (n2746, n_2329, n_2330);
  not g4849 (n_2331, n2745);
  not g4850 (n_2332, n2746);
  and g4851 (n2747, n_2331, n_2332);
  and g4852 (n2748, \a[11] , \a[23] );
  and g4853 (n2749, \a[12] , \a[22] );
  not g4854 (n_2333, n2748);
  not g4855 (n_2334, n2749);
  and g4856 (n2750, n_2333, n_2334);
  and g4857 (n2751, n602, n1919);
  not g4858 (n_2335, n2751);
  not g4861 (n_2336, n2750);
  not g4863 (n_2337, n2754);
  and g4864 (n2755, \a[32] , n_2337);
  and g4865 (n2756, \a[2] , n2755);
  and g4866 (n2757, n_2335, n_2337);
  and g4867 (n2758, n_2336, n2757);
  not g4868 (n_2338, n2756);
  not g4869 (n_2339, n2758);
  and g4870 (n2759, n_2338, n_2339);
  not g4871 (n_2340, n2759);
  and g4872 (n2760, n2747, n_2340);
  not g4873 (n_2341, n2760);
  and g4874 (n2761, n2747, n_2341);
  and g4875 (n2762, n_2340, n_2341);
  not g4876 (n_2342, n2761);
  not g4877 (n_2343, n2762);
  and g4878 (n2763, n_2342, n_2343);
  and g4879 (n2764, n_2296, n_2302);
  and g4880 (n2765, n2763, n2764);
  not g4881 (n_2344, n2763);
  not g4882 (n_2345, n2764);
  and g4883 (n2766, n_2344, n_2345);
  not g4884 (n_2346, n2765);
  not g4885 (n_2347, n2766);
  and g4886 (n2767, n_2346, n_2347);
  and g4887 (n2768, \a[29] , n684);
  and g4888 (n2769, \a[24] , n2768);
  and g4889 (n2770, n484, n1904);
  not g4890 (n_2348, n2769);
  not g4891 (n_2349, n2770);
  and g4892 (n2771, n_2348, n_2349);
  and g4893 (n2772, \a[5] , \a[29] );
  and g4894 (n2773, \a[9] , \a[25] );
  and g4895 (n2774, n2772, n2773);
  not g4896 (n_2350, n2771);
  not g4897 (n_2351, n2774);
  and g4898 (n2775, n_2350, n_2351);
  not g4899 (n_2352, n2775);
  and g4900 (n2776, n_2351, n_2352);
  not g4901 (n_2353, n2772);
  not g4902 (n_2354, n2773);
  and g4903 (n2777, n_2353, n_2354);
  not g4904 (n_2355, n2777);
  and g4905 (n2778, n2776, n_2355);
  and g4906 (n2779, \a[24] , n_2352);
  and g4907 (n2780, \a[10] , n2779);
  not g4908 (n_2356, n2778);
  not g4909 (n_2357, n2780);
  and g4910 (n2781, n_2356, n_2357);
  and g4911 (n2782, n895, n1490);
  and g4912 (n2783, n821, n1492);
  and g4913 (n2784, n745, n1494);
  not g4914 (n_2358, n2783);
  not g4915 (n_2359, n2784);
  and g4916 (n2785, n_2358, n_2359);
  not g4917 (n_2360, n2782);
  not g4918 (n_2361, n2785);
  and g4919 (n2786, n_2360, n_2361);
  not g4920 (n_2362, n2786);
  and g4921 (n2787, \a[21] , n_2362);
  and g4922 (n2788, \a[13] , n2787);
  and g4923 (n2789, n_2360, n_2362);
  and g4924 (n2790, \a[14] , \a[20] );
  and g4925 (n2791, \a[15] , \a[19] );
  not g4926 (n_2363, n2790);
  not g4927 (n_2364, n2791);
  and g4928 (n2792, n_2363, n_2364);
  not g4929 (n_2365, n2792);
  and g4930 (n2793, n2789, n_2365);
  not g4931 (n_2366, n2788);
  not g4932 (n_2367, n2793);
  and g4933 (n2794, n_2366, n_2367);
  not g4934 (n_2368, n2781);
  not g4935 (n_2369, n2794);
  and g4936 (n2795, n_2368, n_2369);
  not g4937 (n_2370, n2795);
  and g4938 (n2796, n_2368, n_2370);
  and g4939 (n2797, n_2369, n_2370);
  not g4940 (n_2371, n2796);
  not g4941 (n_2372, n2797);
  and g4942 (n2798, n_2371, n_2372);
  and g4943 (n2799, n380, n2227);
  and g4944 (n2800, \a[26] , \a[28] );
  and g4945 (n2801, n312, n2800);
  and g4946 (n2802, n335, n2331);
  not g4947 (n_2373, n2801);
  not g4948 (n_2374, n2802);
  and g4949 (n2803, n_2373, n_2374);
  not g4950 (n_2375, n2799);
  not g4951 (n_2376, n2803);
  and g4952 (n2804, n_2375, n_2376);
  not g4953 (n_2377, n2804);
  and g4954 (n2805, \a[28] , n_2377);
  and g4955 (n2806, \a[6] , n2805);
  and g4956 (n2807, n_2375, n_2377);
  and g4957 (n2808, \a[7] , \a[27] );
  and g4958 (n2809, \a[8] , \a[26] );
  not g4959 (n_2378, n2808);
  not g4960 (n_2379, n2809);
  and g4961 (n2810, n_2378, n_2379);
  not g4962 (n_2380, n2810);
  and g4963 (n2811, n2807, n_2380);
  not g4964 (n_2381, n2806);
  not g4965 (n_2382, n2811);
  and g4966 (n2812, n_2381, n_2382);
  not g4967 (n_2383, n2798);
  not g4968 (n_2384, n2812);
  and g4969 (n2813, n_2383, n_2384);
  not g4970 (n_2385, n2813);
  and g4971 (n2814, n_2383, n_2385);
  and g4972 (n2815, n_2384, n_2385);
  not g4973 (n_2386, n2814);
  not g4974 (n_2387, n2815);
  and g4975 (n2816, n_2386, n_2387);
  not g4976 (n_2388, n2816);
  and g4977 (n2817, n2767, n_2388);
  not g4978 (n_2389, n2767);
  and g4979 (n2818, n_2389, n2816);
  and g4980 (n2819, n2604, n2626);
  not g4981 (n_2390, n2604);
  not g4982 (n_2391, n2626);
  and g4983 (n2820, n_2390, n_2391);
  not g4984 (n_2392, n2819);
  not g4985 (n_2393, n2820);
  and g4986 (n2821, n_2392, n_2393);
  not g4987 (n_2394, n2821);
  and g4988 (n2822, n2643, n_2394);
  not g4989 (n_2395, n2643);
  and g4990 (n2823, n_2395, n2821);
  not g4991 (n_2396, n2822);
  not g4992 (n_2397, n2823);
  and g4993 (n2824, n_2396, n_2397);
  and g4994 (n2825, n_2238, n_2250);
  and g4995 (n2826, \a[17] , n2687);
  and g4996 (n2827, \a[1] , \a[33] );
  and g4997 (n2828, n1050, n2827);
  not g4998 (n_2398, n1050);
  not g4999 (n_2399, n2827);
  and g5000 (n2829, n_2398, n_2399);
  not g5001 (n_2400, n2828);
  not g5002 (n_2401, n2829);
  and g5003 (n2830, n_2400, n_2401);
  and g5004 (n2831, n2826, n2830);
  not g5005 (n_2402, n2826);
  not g5006 (n_2403, n2830);
  and g5007 (n2832, n_2402, n_2403);
  not g5008 (n_2404, n2831);
  not g5009 (n_2405, n2832);
  and g5010 (n2833, n_2404, n_2405);
  not g5011 (n_2406, n2658);
  and g5012 (n2834, n_2406, n2833);
  not g5013 (n_2407, n2833);
  and g5014 (n2835, n2658, n_2407);
  not g5015 (n_2408, n2834);
  not g5016 (n_2409, n2835);
  and g5017 (n2836, n_2408, n_2409);
  not g5018 (n_2410, n2825);
  and g5019 (n2837, n_2410, n2836);
  not g5020 (n_2411, n2836);
  and g5021 (n2838, n2825, n_2411);
  not g5022 (n_2412, n2837);
  not g5023 (n_2413, n2838);
  and g5024 (n2839, n_2412, n_2413);
  and g5025 (n2840, n2824, n2839);
  not g5026 (n_2414, n2824);
  not g5027 (n_2415, n2839);
  and g5028 (n2841, n_2414, n_2415);
  not g5029 (n_2416, n2840);
  not g5030 (n_2417, n2841);
  and g5031 (n2842, n_2416, n_2417);
  not g5032 (n_2418, n2818);
  and g5033 (n2843, n_2418, n2842);
  not g5034 (n_2419, n2817);
  and g5035 (n2844, n_2419, n2843);
  not g5036 (n_2420, n2844);
  and g5037 (n2845, n2842, n_2420);
  and g5038 (n2846, n_2418, n_2420);
  and g5039 (n2847, n_2419, n2846);
  not g5040 (n_2421, n2845);
  not g5041 (n_2422, n2847);
  and g5042 (n2848, n_2421, n_2422);
  and g5043 (n2849, n_2306, n_2310);
  and g5044 (n2850, n2848, n2849);
  not g5045 (n_2423, n2848);
  not g5046 (n_2424, n2849);
  and g5047 (n2851, n_2423, n_2424);
  not g5048 (n_2425, n2850);
  not g5049 (n_2426, n2851);
  and g5050 (n2852, n_2425, n_2426);
  and g5051 (n2853, n_2267, n_2271);
  and g5052 (n2854, n2616, n_2254);
  not g5053 (n_2427, n2854);
  and g5054 (n2855, n_2215, n_2427);
  and g5055 (n2856, n_2260, n_2264);
  and g5056 (n2857, n2855, n2856);
  not g5057 (n_2428, n2855);
  not g5058 (n_2429, n2856);
  and g5059 (n2858, n_2428, n_2429);
  not g5060 (n_2430, n2857);
  not g5061 (n_2431, n2858);
  and g5062 (n2859, n_2430, n_2431);
  and g5063 (n2860, n_2196, n_2209);
  and g5064 (n2861, n_2188, n_2192);
  and g5065 (n2862, \a[31] , n202);
  and g5066 (n2863, \a[30] , n212);
  not g5067 (n_2432, n2862);
  not g5068 (n_2433, n2863);
  and g5069 (n2864, n_2432, n_2433);
  and g5070 (n2865, \a[30] , \a[31] );
  and g5071 (n2866, n209, n2865);
  not g5072 (n_2435, n2866);
  and g5073 (n2867, \a[34] , n_2435);
  not g5074 (n_2436, n2864);
  and g5075 (n2868, n_2436, n2867);
  and g5076 (n2869, \a[3] , \a[31] );
  and g5077 (n2870, \a[4] , \a[30] );
  not g5078 (n_2437, n2869);
  not g5079 (n_2438, n2870);
  and g5080 (n2871, n_2437, n_2438);
  not g5081 (n_2439, n2871);
  and g5082 (n2872, n_2435, n_2439);
  and g5083 (n2873, \a[0] , \a[34] );
  not g5084 (n_2440, n2872);
  not g5085 (n_2441, n2873);
  and g5086 (n2874, n_2440, n_2441);
  not g5087 (n_2442, n2868);
  not g5088 (n_2443, n2874);
  and g5089 (n2875, n_2442, n_2443);
  not g5090 (n_2444, n2861);
  and g5091 (n2876, n_2444, n2875);
  not g5092 (n_2445, n2875);
  and g5093 (n2877, n2861, n_2445);
  not g5094 (n_2446, n2876);
  not g5095 (n_2447, n2877);
  and g5096 (n2878, n_2446, n_2447);
  not g5097 (n_2448, n2860);
  and g5098 (n2879, n_2448, n2878);
  not g5099 (n_2449, n2878);
  and g5100 (n2880, n2860, n_2449);
  not g5101 (n_2450, n2879);
  not g5102 (n_2451, n2880);
  and g5103 (n2881, n_2450, n_2451);
  and g5104 (n2882, n2859, n2881);
  not g5105 (n_2452, n2859);
  not g5106 (n_2453, n2881);
  and g5107 (n2883, n_2452, n_2453);
  not g5108 (n_2454, n2882);
  not g5109 (n_2455, n2883);
  and g5110 (n2884, n_2454, n_2455);
  not g5111 (n_2456, n2884);
  and g5112 (n2885, n2853, n_2456);
  not g5113 (n_2457, n2853);
  and g5114 (n2886, n_2457, n2884);
  not g5115 (n_2458, n2885);
  not g5116 (n_2459, n2886);
  and g5117 (n2887, n_2458, n_2459);
  and g5118 (n2888, n2852, n2887);
  not g5119 (n_2460, n2852);
  not g5120 (n_2461, n2887);
  and g5121 (n2889, n_2460, n_2461);
  not g5122 (n_2462, n2888);
  not g5123 (n_2463, n2889);
  and g5124 (n2890, n_2462, n_2463);
  not g5125 (n_2464, n2744);
  and g5126 (n2891, n_2464, n2890);
  not g5127 (n_2465, n2890);
  and g5128 (n2892, n2744, n_2465);
  not g5129 (n_2466, n2891);
  not g5130 (n_2467, n2892);
  and g5131 (n2893, n_2466, n_2467);
  not g5132 (n_2468, n2893);
  and g5133 (n2894, n2743, n_2468);
  not g5134 (n_2469, n2743);
  and g5135 (n2895, n_2469, n_2467);
  and g5136 (n2896, n_2466, n2895);
  not g5137 (n_2470, n2894);
  not g5138 (n_2471, n2896);
  and g5139 (\asquared[35] , n_2470, n_2471);
  not g5140 (n_2472, n2895);
  and g5141 (n2898, n_2466, n_2472);
  and g5142 (n2899, n_2459, n_2462);
  and g5143 (n2900, n_2420, n_2426);
  and g5144 (n2901, n_2393, n_2397);
  and g5145 (n2902, n_2404, n_2408);
  and g5146 (n2903, n2901, n2902);
  not g5147 (n_2473, n2901);
  not g5148 (n_2474, n2902);
  and g5149 (n2904, n_2473, n_2474);
  not g5150 (n_2475, n2903);
  not g5151 (n_2476, n2904);
  and g5152 (n2905, n_2475, n_2476);
  and g5153 (n2906, n_2332, n_2341);
  not g5154 (n_2477, n2905);
  and g5155 (n2907, n_2477, n2906);
  not g5156 (n_2478, n2906);
  and g5157 (n2908, n2905, n_2478);
  not g5158 (n_2479, n2907);
  not g5159 (n_2480, n2908);
  and g5160 (n2909, n_2479, n_2480);
  and g5161 (n2910, n_2412, n_2416);
  not g5162 (n_2481, n2909);
  and g5163 (n2911, n_2481, n2910);
  not g5164 (n_2482, n2910);
  and g5165 (n2912, n2909, n_2482);
  not g5166 (n_2483, n2911);
  not g5167 (n_2484, n2912);
  and g5168 (n2913, n_2483, n_2484);
  and g5169 (n2914, n_2347, n_2419);
  not g5170 (n_2485, n2914);
  and g5171 (n2915, n2913, n_2485);
  not g5172 (n_2486, n2913);
  and g5173 (n2916, n_2486, n2914);
  not g5174 (n_2487, n2915);
  not g5175 (n_2488, n2916);
  and g5176 (n2917, n_2487, n_2488);
  not g5177 (n_2489, n2917);
  and g5178 (n2918, n2900, n_2489);
  not g5179 (n_2490, n2900);
  and g5180 (n2919, n_2490, n2917);
  not g5181 (n_2491, n2918);
  not g5182 (n_2492, n2919);
  and g5183 (n2920, n_2491, n_2492);
  and g5184 (n2921, n312, n2041);
  and g5185 (n2922, \a[27] , \a[30] );
  and g5186 (n2923, n354, n2922);
  and g5187 (n2924, n332, n2617);
  not g5188 (n_2493, n2923);
  not g5189 (n_2494, n2924);
  and g5190 (n2925, n_2493, n_2494);
  not g5191 (n_2495, n2921);
  not g5192 (n_2496, n2925);
  and g5193 (n2926, n_2495, n_2496);
  not g5194 (n_2497, n2926);
  and g5195 (n2927, n_2495, n_2497);
  and g5196 (n2928, \a[6] , \a[29] );
  not g5197 (n_2498, n2229);
  not g5198 (n_2499, n2928);
  and g5199 (n2929, n_2498, n_2499);
  not g5200 (n_2500, n2929);
  and g5201 (n2930, n2927, n_2500);
  and g5202 (n2931, \a[30] , n_2497);
  and g5203 (n2932, \a[5] , n2931);
  not g5204 (n_2501, n2930);
  not g5205 (n_2502, n2932);
  and g5206 (n2933, n_2501, n_2502);
  and g5207 (n2934, \a[16] , \a[19] );
  not g5208 (n_2503, n1052);
  not g5209 (n_2504, n2934);
  and g5210 (n2935, n_2503, n_2504);
  and g5211 (n2936, n1052, n2934);
  not g5212 (n_2505, n2936);
  not g5215 (n_2506, n2935);
  not g5217 (n_2507, n2939);
  and g5218 (n2940, \a[28] , n_2507);
  and g5219 (n2941, \a[7] , n2940);
  and g5220 (n2942, n_2505, n_2507);
  and g5221 (n2943, n_2506, n2942);
  not g5222 (n_2508, n2941);
  not g5223 (n_2509, n2943);
  and g5224 (n2944, n_2508, n_2509);
  not g5225 (n_2510, n2933);
  not g5226 (n_2511, n2944);
  and g5227 (n2945, n_2510, n_2511);
  not g5228 (n_2512, n2945);
  and g5229 (n2946, n_2510, n_2512);
  and g5230 (n2947, n_2511, n_2512);
  not g5231 (n_2513, n2946);
  not g5232 (n_2514, n2947);
  and g5233 (n2948, n_2513, n_2514);
  and g5234 (n2949, \a[9] , \a[26] );
  and g5235 (n2950, \a[10] , \a[25] );
  not g5236 (n_2515, n2949);
  not g5237 (n_2516, n2950);
  and g5238 (n2951, n_2515, n_2516);
  and g5239 (n2952, n484, n2463);
  not g5240 (n_2517, n2952);
  not g5243 (n_2518, n2951);
  not g5245 (n_2519, n2955);
  and g5246 (n2956, \a[31] , n_2519);
  and g5247 (n2957, \a[4] , n2956);
  and g5248 (n2958, n_2517, n_2519);
  and g5249 (n2959, n_2518, n2958);
  not g5250 (n_2520, n2957);
  not g5251 (n_2521, n2959);
  and g5252 (n2960, n_2520, n_2521);
  not g5253 (n_2522, n2948);
  not g5254 (n_2523, n2960);
  and g5255 (n2961, n_2522, n_2523);
  not g5256 (n_2524, n2961);
  and g5257 (n2962, n_2522, n_2524);
  and g5258 (n2963, n_2523, n_2524);
  not g5259 (n_2525, n2962);
  not g5260 (n_2526, n2963);
  and g5261 (n2964, n_2525, n_2526);
  and g5262 (n2965, n_2446, n_2450);
  and g5263 (n2966, n2964, n2965);
  not g5264 (n_2527, n2964);
  not g5265 (n_2528, n2965);
  and g5266 (n2967, n_2527, n_2528);
  not g5267 (n_2529, n2966);
  not g5268 (n_2530, n2967);
  and g5269 (n2968, n_2529, n_2530);
  and g5270 (n2969, \a[0] , \a[35] );
  and g5271 (n2970, \a[2] , \a[33] );
  not g5272 (n_2532, n2969);
  not g5273 (n_2533, n2970);
  and g5274 (n2971, n_2532, n_2533);
  and g5275 (n2972, \a[33] , \a[35] );
  and g5276 (n2973, n196, n2972);
  not g5277 (n_2534, n2971);
  not g5278 (n_2535, n2973);
  and g5279 (n2974, n_2534, n_2535);
  and g5280 (n2975, n2828, n2974);
  not g5281 (n_2536, n2975);
  and g5282 (n2976, n_2535, n_2536);
  and g5283 (n2977, n_2534, n2976);
  and g5284 (n2978, n2828, n_2536);
  not g5285 (n_2537, n2977);
  not g5286 (n_2538, n2978);
  and g5287 (n2979, n_2537, n_2538);
  and g5288 (n2980, \a[3] , \a[32] );
  and g5289 (n2981, \a[11] , \a[24] );
  and g5290 (n2982, \a[12] , \a[23] );
  not g5291 (n_2539, n2981);
  not g5292 (n_2540, n2982);
  and g5293 (n2983, n_2539, n_2540);
  and g5294 (n2984, n602, n1666);
  not g5295 (n_2541, n2984);
  and g5296 (n2985, n2980, n_2541);
  not g5297 (n_2542, n2983);
  and g5298 (n2986, n_2542, n2985);
  not g5299 (n_2543, n2986);
  and g5300 (n2987, n2980, n_2543);
  and g5301 (n2988, n_2541, n_2543);
  and g5302 (n2989, n_2542, n2988);
  not g5303 (n_2544, n2987);
  not g5304 (n_2545, n2989);
  and g5305 (n2990, n_2544, n_2545);
  not g5306 (n_2546, n2979);
  not g5307 (n_2547, n2990);
  and g5308 (n2991, n_2546, n_2547);
  not g5309 (n_2548, n2991);
  and g5310 (n2992, n_2546, n_2548);
  and g5311 (n2993, n_2547, n_2548);
  not g5312 (n_2549, n2992);
  not g5313 (n_2550, n2993);
  and g5314 (n2994, n_2549, n_2550);
  and g5315 (n2995, n895, n1494);
  and g5316 (n2996, n821, n1693);
  and g5317 (n2997, n745, n1574);
  not g5318 (n_2551, n2996);
  not g5319 (n_2552, n2997);
  and g5320 (n2998, n_2551, n_2552);
  not g5321 (n_2553, n2995);
  not g5322 (n_2554, n2998);
  and g5323 (n2999, n_2553, n_2554);
  not g5324 (n_2555, n2999);
  and g5325 (n3000, \a[22] , n_2555);
  and g5326 (n3001, \a[13] , n3000);
  and g5327 (n3002, n_2553, n_2555);
  and g5328 (n3003, \a[14] , \a[21] );
  and g5329 (n3004, \a[15] , \a[20] );
  not g5330 (n_2556, n3003);
  not g5331 (n_2557, n3004);
  and g5332 (n3005, n_2556, n_2557);
  not g5333 (n_2558, n3005);
  and g5334 (n3006, n3002, n_2558);
  not g5335 (n_2559, n3001);
  not g5336 (n_2560, n3006);
  and g5337 (n3007, n_2559, n_2560);
  not g5338 (n_2561, n2994);
  not g5339 (n_2562, n3007);
  and g5340 (n3008, n_2561, n_2562);
  not g5341 (n_2563, n3008);
  and g5342 (n3009, n_2561, n_2563);
  and g5343 (n3010, n_2562, n_2563);
  not g5344 (n_2564, n3009);
  not g5345 (n_2565, n3010);
  and g5346 (n3011, n_2564, n_2565);
  not g5347 (n_2566, n3011);
  and g5348 (n3012, n2968, n_2566);
  not g5349 (n_2567, n2968);
  and g5350 (n3013, n_2567, n3011);
  and g5351 (n3014, n_2431, n_2454);
  and g5352 (n3015, n2757, n2789);
  not g5353 (n_2568, n2757);
  not g5354 (n_2569, n2789);
  and g5355 (n3016, n_2568, n_2569);
  not g5356 (n_2570, n3015);
  not g5357 (n_2571, n3016);
  and g5358 (n3017, n_2570, n_2571);
  and g5359 (n3018, n_2435, n_2442);
  not g5360 (n_2572, n3017);
  and g5361 (n3019, n_2572, n3018);
  not g5362 (n_2573, n3018);
  and g5363 (n3020, n3017, n_2573);
  not g5364 (n_2574, n3019);
  not g5365 (n_2575, n3020);
  and g5366 (n3021, n_2574, n_2575);
  and g5367 (n3022, n_2370, n_2385);
  and g5368 (n3023, \a[34] , n975);
  and g5369 (n3024, \a[1] , \a[34] );
  not g5370 (n_2576, \a[18] );
  not g5371 (n_2577, n3024);
  and g5372 (n3025, n_2576, n_2577);
  not g5373 (n_2578, n3023);
  not g5374 (n_2579, n3025);
  and g5375 (n3026, n_2578, n_2579);
  not g5376 (n_2580, n3026);
  and g5377 (n3027, n2807, n_2580);
  not g5378 (n_2581, n2807);
  and g5379 (n3028, n_2581, n3026);
  not g5380 (n_2582, n3027);
  not g5381 (n_2583, n3028);
  and g5382 (n3029, n_2582, n_2583);
  not g5383 (n_2584, n2776);
  and g5384 (n3030, n_2584, n3029);
  not g5385 (n_2585, n3029);
  and g5386 (n3031, n2776, n_2585);
  not g5387 (n_2586, n3030);
  not g5388 (n_2587, n3031);
  and g5389 (n3032, n_2586, n_2587);
  not g5390 (n_2588, n3022);
  and g5391 (n3033, n_2588, n3032);
  not g5392 (n_2589, n3032);
  and g5393 (n3034, n3022, n_2589);
  not g5394 (n_2590, n3033);
  not g5395 (n_2591, n3034);
  and g5396 (n3035, n_2590, n_2591);
  and g5397 (n3036, n3021, n3035);
  not g5398 (n_2592, n3021);
  not g5399 (n_2593, n3035);
  and g5400 (n3037, n_2592, n_2593);
  not g5401 (n_2594, n3036);
  not g5402 (n_2595, n3037);
  and g5403 (n3038, n_2594, n_2595);
  not g5404 (n_2596, n3014);
  and g5405 (n3039, n_2596, n3038);
  not g5406 (n_2597, n3038);
  and g5407 (n3040, n3014, n_2597);
  not g5408 (n_2598, n3039);
  not g5409 (n_2599, n3040);
  and g5410 (n3041, n_2598, n_2599);
  not g5411 (n_2600, n3013);
  and g5412 (n3042, n_2600, n3041);
  not g5413 (n_2601, n3012);
  and g5414 (n3043, n_2601, n3042);
  not g5415 (n_2602, n3043);
  and g5416 (n3044, n3041, n_2602);
  and g5417 (n3045, n_2600, n_2602);
  and g5418 (n3046, n_2601, n3045);
  not g5419 (n_2603, n3044);
  not g5420 (n_2604, n3046);
  and g5421 (n3047, n_2603, n_2604);
  not g5422 (n_2605, n2920);
  and g5423 (n3048, n_2605, n3047);
  not g5424 (n_2606, n3047);
  and g5425 (n3049, n2920, n_2606);
  not g5426 (n_2607, n3048);
  not g5427 (n_2608, n3049);
  and g5428 (n3050, n_2607, n_2608);
  not g5429 (n_2609, n3050);
  and g5430 (n3051, n2899, n_2609);
  not g5431 (n_2610, n2899);
  and g5432 (n3052, n_2610, n3050);
  not g5433 (n_2611, n3051);
  not g5434 (n_2612, n3052);
  and g5435 (n3053, n_2611, n_2612);
  not g5436 (n_2613, n2898);
  not g5437 (n_2614, n3053);
  and g5438 (n3054, n_2613, n_2614);
  and g5439 (n3055, n2898, n3053);
  or g5440 (\asquared[36] , n3054, n3055);
  and g5441 (n3057, n_2492, n_2608);
  and g5442 (n3058, n_2598, n_2602);
  and g5443 (n3059, n_2571, n_2575);
  and g5444 (n3060, n_2583, n_2586);
  and g5445 (n3061, n3059, n3060);
  not g5446 (n_2615, n3059);
  not g5447 (n_2616, n3060);
  and g5448 (n3062, n_2615, n_2616);
  not g5449 (n_2617, n3061);
  not g5450 (n_2618, n3062);
  and g5451 (n3063, n_2617, n_2618);
  and g5452 (n3064, n_2548, n_2563);
  not g5453 (n_2619, n3063);
  and g5454 (n3065, n_2619, n3064);
  not g5455 (n_2620, n3064);
  and g5456 (n3066, n3063, n_2620);
  not g5457 (n_2621, n3065);
  not g5458 (n_2622, n3066);
  and g5459 (n3067, n_2621, n_2622);
  and g5460 (n3068, n_2590, n_2594);
  not g5461 (n_2623, n3067);
  and g5462 (n3069, n_2623, n3068);
  not g5463 (n_2624, n3068);
  and g5464 (n3070, n3067, n_2624);
  not g5465 (n_2625, n3069);
  not g5466 (n_2626, n3070);
  and g5467 (n3071, n_2625, n_2626);
  and g5468 (n3072, n_2530, n_2601);
  not g5469 (n_2627, n3072);
  and g5470 (n3073, n3071, n_2627);
  not g5471 (n_2628, n3071);
  and g5472 (n3074, n_2628, n3072);
  not g5473 (n_2629, n3073);
  not g5474 (n_2630, n3074);
  and g5475 (n3075, n_2629, n_2630);
  not g5476 (n_2631, n3058);
  and g5477 (n3076, n_2631, n3075);
  not g5478 (n_2632, n3075);
  and g5479 (n3077, n3058, n_2632);
  not g5480 (n_2633, n3076);
  not g5481 (n_2634, n3077);
  and g5482 (n3078, n_2633, n_2634);
  and g5483 (n3079, \a[12] , \a[24] );
  and g5484 (n3080, \a[13] , \a[23] );
  not g5485 (n_2635, n3079);
  not g5486 (n_2636, n3080);
  and g5487 (n3081, n_2635, n_2636);
  and g5488 (n3082, n748, n1666);
  not g5489 (n_2637, n3082);
  not g5492 (n_2638, n3081);
  not g5494 (n_2639, n3085);
  and g5495 (n3086, n_2637, n_2639);
  and g5496 (n3087, n_2638, n3086);
  and g5497 (n3088, \a[34] , n_2639);
  and g5498 (n3089, \a[2] , n3088);
  not g5499 (n_2640, n3087);
  not g5500 (n_2641, n3089);
  and g5501 (n3090, n_2640, n_2641);
  and g5502 (n3091, \a[9] , \a[31] );
  and g5503 (n3092, n2451, n3091);
  and g5504 (n3093, n484, n2227);
  and g5505 (n3094, n2309, n2352);
  not g5506 (n_2642, n3093);
  not g5507 (n_2643, n3094);
  and g5508 (n3095, n_2642, n_2643);
  not g5509 (n_2644, n3092);
  not g5510 (n_2645, n3095);
  and g5511 (n3096, n_2644, n_2645);
  not g5512 (n_2646, n3096);
  and g5513 (n3097, \a[26] , n_2646);
  and g5514 (n3098, \a[10] , n3097);
  and g5515 (n3099, n_2644, n_2646);
  and g5516 (n3100, \a[5] , \a[31] );
  and g5517 (n3101, \a[9] , \a[27] );
  not g5518 (n_2647, n3100);
  not g5519 (n_2648, n3101);
  and g5520 (n3102, n_2647, n_2648);
  not g5521 (n_2649, n3102);
  and g5522 (n3103, n3099, n_2649);
  not g5523 (n_2650, n3098);
  not g5524 (n_2651, n3103);
  and g5525 (n3104, n_2650, n_2651);
  not g5526 (n_2652, n3090);
  not g5527 (n_2653, n3104);
  and g5528 (n3105, n_2652, n_2653);
  not g5529 (n_2654, n3105);
  and g5530 (n3106, n_2652, n_2654);
  and g5531 (n3107, n_2653, n_2654);
  not g5532 (n_2655, n3106);
  not g5533 (n_2656, n3107);
  and g5534 (n3108, n_2655, n_2656);
  and g5535 (n3109, n380, n2334);
  and g5536 (n3110, \a[28] , \a[30] );
  and g5537 (n3111, n312, n3110);
  and g5538 (n3112, n335, n2617);
  not g5539 (n_2657, n3111);
  not g5540 (n_2658, n3112);
  and g5541 (n3113, n_2657, n_2658);
  not g5542 (n_2659, n3109);
  not g5543 (n_2660, n3113);
  and g5544 (n3114, n_2659, n_2660);
  not g5545 (n_2661, n3114);
  and g5546 (n3115, \a[30] , n_2661);
  and g5547 (n3116, \a[6] , n3115);
  and g5548 (n3117, n_2659, n_2661);
  and g5549 (n3118, \a[7] , \a[29] );
  and g5550 (n3119, \a[8] , \a[28] );
  not g5551 (n_2662, n3118);
  not g5552 (n_2663, n3119);
  and g5553 (n3120, n_2662, n_2663);
  not g5554 (n_2664, n3120);
  and g5555 (n3121, n3117, n_2664);
  not g5556 (n_2665, n3116);
  not g5557 (n_2666, n3121);
  and g5558 (n3122, n_2665, n_2666);
  not g5559 (n_2667, n3108);
  not g5560 (n_2668, n3122);
  and g5561 (n3123, n_2667, n_2668);
  not g5562 (n_2669, n3123);
  and g5563 (n3124, n_2667, n_2669);
  and g5564 (n3125, n_2668, n_2669);
  not g5565 (n_2670, n3124);
  not g5566 (n_2671, n3125);
  and g5567 (n3126, n_2670, n_2671);
  and g5568 (n3127, n_2476, n_2480);
  and g5569 (n3128, \a[0] , \a[36] );
  and g5570 (n3129, n3023, n3128);
  not g5571 (n_2673, n3129);
  and g5572 (n3130, n3023, n_2673);
  and g5573 (n3131, n_2578, n3128);
  not g5574 (n_2674, n3130);
  not g5575 (n_2675, n3131);
  and g5576 (n3132, n_2674, n_2675);
  and g5577 (n3133, \a[1] , \a[35] );
  and g5578 (n3134, \a[17] , \a[19] );
  and g5579 (n3135, n3133, n3134);
  not g5580 (n_2676, n3135);
  and g5581 (n3136, n3133, n_2676);
  and g5582 (n3137, n3134, n_2676);
  not g5583 (n_2677, n3136);
  not g5584 (n_2678, n3137);
  and g5585 (n3138, n_2677, n_2678);
  not g5586 (n_2679, n3132);
  not g5587 (n_2680, n3138);
  and g5588 (n3139, n_2679, n_2680);
  not g5589 (n_2681, n3139);
  and g5590 (n3140, n_2679, n_2681);
  and g5591 (n3141, n_2680, n_2681);
  not g5592 (n_2682, n3140);
  not g5593 (n_2683, n3141);
  and g5594 (n3142, n_2682, n_2683);
  and g5595 (n3143, \a[32] , \a[33] );
  and g5596 (n3144, n209, n3143);
  and g5597 (n3145, \a[11] , \a[25] );
  and g5598 (n3146, \a[3] , \a[33] );
  and g5599 (n3147, n3145, n3146);
  not g5600 (n_2684, n3144);
  not g5601 (n_2685, n3147);
  and g5602 (n3148, n_2684, n_2685);
  and g5603 (n3149, \a[4] , \a[32] );
  and g5604 (n3150, n3145, n3149);
  not g5605 (n_2686, n3148);
  not g5606 (n_2687, n3150);
  and g5607 (n3151, n_2686, n_2687);
  not g5608 (n_2688, n3151);
  and g5609 (n3152, n_2687, n_2688);
  not g5610 (n_2689, n3145);
  not g5611 (n_2690, n3149);
  and g5612 (n3153, n_2689, n_2690);
  not g5613 (n_2691, n3153);
  and g5614 (n3154, n3152, n_2691);
  and g5615 (n3155, n3146, n_2688);
  not g5616 (n_2692, n3154);
  not g5617 (n_2693, n3155);
  and g5618 (n3156, n_2692, n_2693);
  and g5619 (n3157, n891, n1494);
  and g5620 (n3158, n893, n1693);
  and g5621 (n3159, n895, n1574);
  not g5622 (n_2694, n3158);
  not g5623 (n_2695, n3159);
  and g5624 (n3160, n_2694, n_2695);
  not g5625 (n_2696, n3157);
  not g5626 (n_2697, n3160);
  and g5627 (n3161, n_2696, n_2697);
  not g5628 (n_2698, n3161);
  and g5629 (n3162, \a[22] , n_2698);
  and g5630 (n3163, \a[14] , n3162);
  and g5631 (n3164, n_2696, n_2698);
  and g5632 (n3165, \a[15] , \a[21] );
  and g5633 (n3166, \a[16] , \a[20] );
  not g5634 (n_2699, n3165);
  not g5635 (n_2700, n3166);
  and g5636 (n3167, n_2699, n_2700);
  not g5637 (n_2701, n3167);
  and g5638 (n3168, n3164, n_2701);
  not g5639 (n_2702, n3163);
  not g5640 (n_2703, n3168);
  and g5641 (n3169, n_2702, n_2703);
  not g5642 (n_2704, n3156);
  not g5643 (n_2705, n3169);
  and g5644 (n3170, n_2704, n_2705);
  not g5645 (n_2706, n3170);
  and g5646 (n3171, n_2704, n_2706);
  and g5647 (n3172, n_2705, n_2706);
  not g5648 (n_2707, n3171);
  not g5649 (n_2708, n3172);
  and g5650 (n3173, n_2707, n_2708);
  not g5651 (n_2709, n3142);
  and g5652 (n3174, n_2709, n3173);
  not g5653 (n_2710, n3173);
  and g5654 (n3175, n3142, n_2710);
  not g5655 (n_2711, n3174);
  not g5656 (n_2712, n3175);
  and g5657 (n3176, n_2711, n_2712);
  not g5658 (n_2713, n3127);
  not g5659 (n_2714, n3176);
  and g5660 (n3177, n_2713, n_2714);
  not g5661 (n_2715, n3177);
  and g5662 (n3178, n_2713, n_2715);
  and g5663 (n3179, n_2714, n_2715);
  not g5664 (n_2716, n3178);
  not g5665 (n_2717, n3179);
  and g5666 (n3180, n_2716, n_2717);
  not g5667 (n_2718, n3126);
  not g5668 (n_2719, n3180);
  and g5669 (n3181, n_2718, n_2719);
  not g5670 (n_2720, n3181);
  and g5671 (n3182, n_2718, n_2720);
  and g5672 (n3183, n_2719, n_2720);
  not g5673 (n_2721, n3182);
  not g5674 (n_2722, n3183);
  and g5675 (n3184, n_2721, n_2722);
  and g5676 (n3185, n_2484, n_2487);
  and g5677 (n3186, n2927, n2958);
  not g5678 (n_2723, n2927);
  not g5679 (n_2724, n2958);
  and g5680 (n3187, n_2723, n_2724);
  not g5681 (n_2725, n3186);
  not g5682 (n_2726, n3187);
  and g5683 (n3188, n_2725, n_2726);
  not g5684 (n_2727, n3188);
  and g5685 (n3189, n2942, n_2727);
  not g5686 (n_2728, n2942);
  and g5687 (n3190, n_2728, n3188);
  not g5688 (n_2729, n3189);
  not g5689 (n_2730, n3190);
  and g5690 (n3191, n_2729, n_2730);
  and g5691 (n3192, n2988, n3002);
  not g5692 (n_2731, n2988);
  not g5693 (n_2732, n3002);
  and g5694 (n3193, n_2731, n_2732);
  not g5695 (n_2733, n3192);
  not g5696 (n_2734, n3193);
  and g5697 (n3194, n_2733, n_2734);
  not g5698 (n_2735, n3194);
  and g5699 (n3195, n2976, n_2735);
  not g5700 (n_2736, n2976);
  and g5701 (n3196, n_2736, n3194);
  not g5702 (n_2737, n3195);
  not g5703 (n_2738, n3196);
  and g5704 (n3197, n_2737, n_2738);
  and g5705 (n3198, n_2512, n_2524);
  not g5706 (n_2739, n3197);
  and g5707 (n3199, n_2739, n3198);
  not g5708 (n_2740, n3198);
  and g5709 (n3200, n3197, n_2740);
  not g5710 (n_2741, n3199);
  not g5711 (n_2742, n3200);
  and g5712 (n3201, n_2741, n_2742);
  and g5713 (n3202, n3191, n3201);
  not g5714 (n_2743, n3191);
  not g5715 (n_2744, n3201);
  and g5716 (n3203, n_2743, n_2744);
  not g5717 (n_2745, n3202);
  not g5718 (n_2746, n3203);
  and g5719 (n3204, n_2745, n_2746);
  not g5720 (n_2747, n3185);
  and g5721 (n3205, n_2747, n3204);
  not g5722 (n_2748, n3205);
  and g5723 (n3206, n_2747, n_2748);
  and g5724 (n3207, n3204, n_2748);
  not g5725 (n_2749, n3206);
  not g5726 (n_2750, n3207);
  and g5727 (n3208, n_2749, n_2750);
  not g5728 (n_2751, n3184);
  not g5729 (n_2752, n3208);
  and g5730 (n3209, n_2751, n_2752);
  and g5731 (n3210, n3184, n_2750);
  and g5732 (n3211, n_2749, n3210);
  not g5733 (n_2753, n3209);
  not g5734 (n_2754, n3211);
  and g5735 (n3212, n_2753, n_2754);
  and g5736 (n3213, n3078, n3212);
  not g5737 (n_2755, n3078);
  not g5738 (n_2756, n3212);
  and g5739 (n3214, n_2755, n_2756);
  not g5740 (n_2757, n3213);
  not g5741 (n_2758, n3214);
  and g5742 (n3215, n_2757, n_2758);
  not g5743 (n_2759, n3215);
  and g5744 (n3216, n3057, n_2759);
  not g5745 (n_2760, n3057);
  and g5746 (n3217, n_2760, n3215);
  not g5747 (n_2761, n3216);
  not g5748 (n_2762, n3217);
  and g5749 (n3218, n_2761, n_2762);
  and g5750 (n3219, n_2613, n_2611);
  not g5751 (n_2763, n3219);
  and g5752 (n3220, n_2612, n_2763);
  not g5753 (n_2764, n3218);
  and g5754 (n3221, n_2764, n3220);
  not g5755 (n_2765, n3220);
  and g5756 (n3222, n3218, n_2765);
  not g5757 (n_2766, n3221);
  not g5758 (n_2767, n3222);
  and g5759 (\asquared[37] , n_2766, n_2767);
  and g5760 (n3224, n_2633, n_2757);
  and g5761 (n3225, n_2626, n_2629);
  and g5762 (n3226, n_2673, n_2681);
  and g5763 (n3227, n3099, n3226);
  not g5764 (n_2768, n3099);
  not g5765 (n_2769, n3226);
  and g5766 (n3228, n_2768, n_2769);
  not g5767 (n_2770, n3227);
  not g5768 (n_2771, n3228);
  and g5769 (n3229, n_2770, n_2771);
  and g5770 (n3230, n895, n1919);
  and g5771 (n3231, n821, n2115);
  and g5772 (n3232, n745, n1666);
  not g5773 (n_2772, n3231);
  not g5774 (n_2773, n3232);
  and g5775 (n3233, n_2772, n_2773);
  not g5776 (n_2774, n3230);
  not g5777 (n_2775, n3233);
  and g5778 (n3234, n_2774, n_2775);
  not g5779 (n_2776, n3234);
  and g5780 (n3235, \a[24] , n_2776);
  and g5781 (n3236, \a[13] , n3235);
  and g5782 (n3237, \a[14] , \a[23] );
  and g5783 (n3238, \a[15] , \a[22] );
  not g5784 (n_2777, n3237);
  not g5785 (n_2778, n3238);
  and g5786 (n3239, n_2777, n_2778);
  and g5787 (n3240, n_2774, n_2776);
  not g5788 (n_2779, n3239);
  and g5789 (n3241, n_2779, n3240);
  not g5790 (n_2780, n3236);
  not g5791 (n_2781, n3241);
  and g5792 (n3242, n_2780, n_2781);
  not g5793 (n_2782, n3242);
  and g5794 (n3243, n3229, n_2782);
  not g5795 (n_2783, n3243);
  and g5796 (n3244, n3229, n_2783);
  and g5797 (n3245, n_2782, n_2783);
  not g5798 (n_2784, n3244);
  not g5799 (n_2785, n3245);
  and g5800 (n3246, n_2784, n_2785);
  and g5801 (n3247, n3152, n3164);
  not g5802 (n_2786, n3152);
  not g5803 (n_2787, n3164);
  and g5804 (n3248, n_2786, n_2787);
  not g5805 (n_2788, n3247);
  not g5806 (n_2789, n3248);
  and g5807 (n3249, n_2788, n_2789);
  not g5808 (n_2790, n3249);
  and g5809 (n3250, n3086, n_2790);
  not g5810 (n_2791, n3086);
  and g5811 (n3251, n_2791, n3249);
  not g5812 (n_2792, n3250);
  not g5813 (n_2793, n3251);
  and g5814 (n3252, n_2792, n_2793);
  and g5815 (n3253, n_2709, n_2710);
  not g5816 (n_2794, n3253);
  and g5817 (n3254, n_2706, n_2794);
  not g5818 (n_2795, n3254);
  and g5819 (n3255, n3252, n_2795);
  not g5820 (n_2796, n3252);
  and g5821 (n3256, n_2796, n3254);
  not g5822 (n_2797, n3255);
  not g5823 (n_2798, n3256);
  and g5824 (n3257, n_2797, n_2798);
  and g5825 (n3258, n3246, n3257);
  not g5826 (n_2799, n3246);
  not g5827 (n_2800, n3257);
  and g5828 (n3259, n_2799, n_2800);
  not g5829 (n_2801, n3258);
  not g5830 (n_2802, n3259);
  and g5831 (n3260, n_2801, n_2802);
  not g5832 (n_2803, n3225);
  not g5833 (n_2804, n3260);
  and g5834 (n3261, n_2803, n_2804);
  and g5835 (n3262, n3225, n3260);
  not g5836 (n_2805, n3261);
  not g5837 (n_2806, n3262);
  and g5838 (n3263, n_2805, n_2806);
  and g5839 (n3264, \a[10] , \a[32] );
  and g5840 (n3265, n2451, n3264);
  and g5841 (n3266, \a[26] , \a[32] );
  and g5842 (n3267, n502, n3266);
  and g5843 (n3268, n723, n2227);
  not g5844 (n_2807, n3267);
  not g5845 (n_2808, n3268);
  and g5846 (n3269, n_2807, n_2808);
  not g5847 (n_2809, n3265);
  not g5848 (n_2810, n3269);
  and g5849 (n3270, n_2809, n_2810);
  not g5850 (n_2811, n3270);
  and g5851 (n3271, n_2809, n_2811);
  and g5852 (n3272, \a[5] , \a[32] );
  and g5853 (n3273, \a[10] , \a[27] );
  not g5854 (n_2812, n3272);
  not g5855 (n_2813, n3273);
  and g5856 (n3274, n_2812, n_2813);
  not g5857 (n_2814, n3274);
  and g5858 (n3275, n3271, n_2814);
  and g5859 (n3276, \a[26] , n_2811);
  and g5860 (n3277, \a[11] , n3276);
  not g5861 (n_2815, n3275);
  not g5862 (n_2816, n3277);
  and g5863 (n3278, n_2815, n_2816);
  not g5864 (n_2817, n1149);
  not g5865 (n_2818, n1333);
  and g5866 (n3279, n_2817, n_2818);
  and g5867 (n3280, n1052, n1490);
  not g5868 (n_2819, n3280);
  not g5871 (n_2820, n3279);
  not g5873 (n_2821, n3283);
  and g5874 (n3284, \a[29] , n_2821);
  and g5875 (n3285, \a[8] , n3284);
  and g5876 (n3286, n_2819, n_2821);
  and g5877 (n3287, n_2820, n3286);
  not g5878 (n_2822, n3285);
  not g5879 (n_2823, n3287);
  and g5880 (n3288, n_2822, n_2823);
  not g5881 (n_2824, n3278);
  not g5882 (n_2825, n3288);
  and g5883 (n3289, n_2824, n_2825);
  not g5884 (n_2826, n3289);
  and g5885 (n3290, n_2824, n_2826);
  and g5886 (n3291, n_2825, n_2826);
  not g5887 (n_2827, n3290);
  not g5888 (n_2828, n3291);
  and g5889 (n3292, n_2827, n_2828);
  and g5890 (n3293, n_2734, n_2738);
  and g5891 (n3294, n3292, n3293);
  not g5892 (n_2829, n3292);
  not g5893 (n_2830, n3293);
  and g5894 (n3295, n_2829, n_2830);
  not g5895 (n_2831, n3294);
  not g5896 (n_2832, n3295);
  and g5897 (n3296, n_2831, n_2832);
  and g5898 (n3297, n_2618, n_2622);
  not g5899 (n_2833, n3296);
  and g5900 (n3298, n_2833, n3297);
  not g5901 (n_2834, n3297);
  and g5902 (n3299, n3296, n_2834);
  not g5903 (n_2835, n3298);
  not g5904 (n_2836, n3299);
  and g5905 (n3300, n_2835, n_2836);
  and g5906 (n3301, \a[25] , \a[33] );
  and g5907 (n3302, n744, n3301);
  and g5908 (n3303, \a[25] , n482);
  and g5909 (n3304, \a[33] , n212);
  not g5910 (n_2837, n3303);
  not g5911 (n_2838, n3304);
  and g5912 (n3305, n_2837, n_2838);
  not g5913 (n_2840, n3302);
  and g5914 (n3306, \a[37] , n_2840);
  not g5915 (n_2841, n3305);
  and g5916 (n3307, n_2841, n3306);
  not g5917 (n_2842, n3307);
  and g5918 (n3308, n_2840, n_2842);
  and g5919 (n3309, \a[4] , \a[33] );
  and g5920 (n3310, \a[12] , \a[25] );
  not g5921 (n_2843, n3309);
  not g5922 (n_2844, n3310);
  and g5923 (n3311, n_2843, n_2844);
  not g5924 (n_2845, n3311);
  and g5925 (n3312, n3308, n_2845);
  and g5926 (n3313, \a[37] , n_2842);
  and g5927 (n3314, \a[0] , n3313);
  not g5928 (n_2846, n3312);
  not g5929 (n_2847, n3314);
  and g5930 (n3315, n_2846, n_2847);
  and g5931 (n3316, \a[2] , \a[35] );
  and g5932 (n3317, \a[3] , \a[34] );
  not g5933 (n_2848, n3316);
  not g5934 (n_2849, n3317);
  and g5935 (n3318, n_2848, n_2849);
  and g5936 (n3319, \a[34] , \a[35] );
  and g5937 (n3320, n218, n3319);
  not g5938 (n_2850, n3320);
  not g5941 (n_2851, n3318);
  not g5943 (n_2852, n3323);
  and g5944 (n3324, \a[21] , n_2852);
  and g5945 (n3325, \a[16] , n3324);
  and g5946 (n3326, n_2850, n_2852);
  and g5947 (n3327, n_2851, n3326);
  not g5948 (n_2853, n3325);
  not g5949 (n_2854, n3327);
  and g5950 (n3328, n_2853, n_2854);
  not g5951 (n_2855, n3315);
  not g5952 (n_2856, n3328);
  and g5953 (n3329, n_2855, n_2856);
  not g5954 (n_2857, n3329);
  and g5955 (n3330, n_2855, n_2857);
  and g5956 (n3331, n_2856, n_2857);
  not g5957 (n_2858, n3330);
  not g5958 (n_2859, n3331);
  and g5959 (n3332, n_2858, n_2859);
  and g5960 (n3333, \a[9] , \a[28] );
  and g5961 (n3334, n335, n2865);
  and g5962 (n3335, n763, n3110);
  and g5963 (n3336, \a[6] , \a[31] );
  and g5964 (n3337, n3333, n3336);
  not g5965 (n_2860, n3335);
  not g5966 (n_2861, n3337);
  and g5967 (n3338, n_2860, n_2861);
  not g5968 (n_2862, n3334);
  not g5969 (n_2863, n3338);
  and g5970 (n3339, n_2862, n_2863);
  not g5971 (n_2864, n3339);
  and g5972 (n3340, n3333, n_2864);
  and g5973 (n3341, n_2862, n_2864);
  and g5974 (n3342, \a[7] , \a[30] );
  not g5975 (n_2865, n3336);
  not g5976 (n_2866, n3342);
  and g5977 (n3343, n_2865, n_2866);
  not g5978 (n_2867, n3343);
  and g5979 (n3344, n3341, n_2867);
  not g5980 (n_2868, n3340);
  not g5981 (n_2869, n3344);
  and g5982 (n3345, n_2868, n_2869);
  not g5983 (n_2870, n3332);
  not g5984 (n_2871, n3345);
  and g5985 (n3346, n_2870, n_2871);
  not g5986 (n_2872, n3346);
  and g5987 (n3347, n_2870, n_2872);
  and g5988 (n3348, n_2871, n_2872);
  not g5989 (n_2873, n3347);
  not g5990 (n_2874, n3348);
  and g5991 (n3349, n_2873, n_2874);
  not g5992 (n_2875, n3300);
  and g5993 (n3350, n_2875, n3349);
  not g5994 (n_2876, n3349);
  and g5995 (n3351, n3300, n_2876);
  not g5996 (n_2877, n3350);
  not g5997 (n_2878, n3351);
  and g5998 (n3352, n_2877, n_2878);
  and g5999 (n3353, n3263, n3352);
  not g6000 (n_2879, n3263);
  not g6001 (n_2880, n3352);
  and g6002 (n3354, n_2879, n_2880);
  not g6003 (n_2881, n3353);
  not g6004 (n_2882, n3354);
  and g6005 (n3355, n_2881, n_2882);
  and g6006 (n3356, n_2748, n_2753);
  and g6007 (n3357, n_2715, n_2720);
  and g6008 (n3358, n_2742, n_2745);
  and g6009 (n3359, n_2654, n_2669);
  and g6010 (n3360, n_2726, n_2730);
  and g6011 (n3361, \a[36] , n1077);
  and g6012 (n3362, \a[1] , \a[36] );
  not g6013 (n_2883, \a[19] );
  not g6014 (n_2884, n3362);
  and g6015 (n3363, n_2883, n_2884);
  not g6016 (n_2885, n3361);
  not g6017 (n_2886, n3363);
  and g6018 (n3364, n_2885, n_2886);
  and g6019 (n3365, n3135, n3364);
  not g6020 (n_2887, n3365);
  and g6021 (n3366, n3135, n_2887);
  and g6022 (n3367, n3364, n_2887);
  not g6023 (n_2888, n3366);
  not g6024 (n_2889, n3367);
  and g6025 (n3368, n_2888, n_2889);
  not g6026 (n_2890, n3117);
  not g6027 (n_2891, n3368);
  and g6028 (n3369, n_2890, n_2891);
  and g6029 (n3370, n3117, n_2889);
  and g6030 (n3371, n_2888, n3370);
  not g6031 (n_2892, n3369);
  not g6032 (n_2893, n3371);
  and g6033 (n3372, n_2892, n_2893);
  not g6034 (n_2894, n3360);
  and g6035 (n3373, n_2894, n3372);
  not g6036 (n_2895, n3372);
  and g6037 (n3374, n3360, n_2895);
  not g6038 (n_2896, n3373);
  not g6039 (n_2897, n3374);
  and g6040 (n3375, n_2896, n_2897);
  not g6041 (n_2898, n3359);
  and g6042 (n3376, n_2898, n3375);
  not g6043 (n_2899, n3375);
  and g6044 (n3377, n3359, n_2899);
  not g6045 (n_2900, n3376);
  not g6046 (n_2901, n3377);
  and g6047 (n3378, n_2900, n_2901);
  not g6048 (n_2902, n3358);
  and g6049 (n3379, n_2902, n3378);
  not g6050 (n_2903, n3378);
  and g6051 (n3380, n3358, n_2903);
  not g6052 (n_2904, n3379);
  not g6053 (n_2905, n3380);
  and g6054 (n3381, n_2904, n_2905);
  not g6055 (n_2906, n3357);
  and g6056 (n3382, n_2906, n3381);
  not g6057 (n_2907, n3381);
  and g6058 (n3383, n3357, n_2907);
  not g6059 (n_2908, n3382);
  not g6060 (n_2909, n3383);
  and g6061 (n3384, n_2908, n_2909);
  not g6062 (n_2910, n3356);
  and g6063 (n3385, n_2910, n3384);
  not g6064 (n_2911, n3385);
  and g6065 (n3386, n_2910, n_2911);
  and g6066 (n3387, n3384, n_2911);
  not g6067 (n_2912, n3386);
  not g6068 (n_2913, n3387);
  and g6069 (n3388, n_2912, n_2913);
  not g6070 (n_2914, n3388);
  and g6071 (n3389, n3355, n_2914);
  not g6072 (n_2915, n3355);
  and g6073 (n3390, n_2915, n_2913);
  and g6074 (n3391, n_2912, n3390);
  not g6075 (n_2916, n3389);
  not g6076 (n_2917, n3391);
  and g6077 (n3392, n_2916, n_2917);
  not g6078 (n_2918, n3224);
  and g6079 (n3393, n_2918, n3392);
  not g6080 (n_2919, n3392);
  and g6081 (n3394, n3224, n_2919);
  not g6082 (n_2920, n3393);
  not g6083 (n_2921, n3394);
  and g6084 (n3395, n_2920, n_2921);
  and g6085 (n3396, n_2761, n_2765);
  not g6086 (n_2922, n3396);
  and g6087 (n3397, n_2762, n_2922);
  not g6088 (n_2923, n3395);
  and g6089 (n3398, n_2923, n3397);
  not g6090 (n_2924, n3397);
  and g6091 (n3399, n3395, n_2924);
  not g6092 (n_2925, n3398);
  not g6093 (n_2926, n3399);
  and g6094 (\asquared[38] , n_2925, n_2926);
  and g6095 (n3401, n_2911, n_2916);
  and g6096 (n3402, n_2836, n_2878);
  and g6097 (n3403, n_2799, n3257);
  not g6098 (n_2927, n3403);
  and g6099 (n3404, n_2797, n_2927);
  not g6100 (n_2928, n3402);
  not g6101 (n_2929, n3404);
  and g6102 (n3405, n_2928, n_2929);
  not g6103 (n_2930, n3405);
  and g6104 (n3406, n_2928, n_2930);
  and g6105 (n3407, n_2929, n_2930);
  not g6106 (n_2931, n3406);
  not g6107 (n_2932, n3407);
  and g6108 (n3408, n_2931, n_2932);
  and g6109 (n3409, n3308, n3326);
  not g6110 (n_2933, n3308);
  not g6111 (n_2934, n3326);
  and g6112 (n3410, n_2933, n_2934);
  not g6113 (n_2935, n3409);
  not g6114 (n_2936, n3410);
  and g6115 (n3411, n_2935, n_2936);
  not g6116 (n_2937, n3411);
  and g6117 (n3412, n3240, n_2937);
  not g6118 (n_2938, n3240);
  and g6119 (n3413, n_2938, n3411);
  not g6120 (n_2939, n3412);
  not g6121 (n_2940, n3413);
  and g6122 (n3414, n_2939, n_2940);
  and g6123 (n3415, n_2826, n_2832);
  not g6124 (n_2941, n3414);
  and g6125 (n3416, n_2941, n3415);
  not g6126 (n_2942, n3415);
  and g6127 (n3417, n3414, n_2942);
  not g6128 (n_2943, n3416);
  not g6129 (n_2944, n3417);
  and g6130 (n3418, n_2943, n_2944);
  and g6131 (n3419, \a[6] , \a[32] );
  and g6132 (n3420, \a[10] , \a[28] );
  not g6133 (n_2945, n3419);
  not g6134 (n_2946, n3420);
  and g6135 (n3421, n_2945, n_2946);
  and g6136 (n3422, n332, n3143);
  and g6137 (n3423, \a[5] , \a[33] );
  and g6138 (n3424, n3420, n3423);
  not g6139 (n_2947, n3422);
  not g6140 (n_2948, n3424);
  and g6141 (n3425, n_2947, n_2948);
  and g6142 (n3426, n3419, n3420);
  not g6143 (n_2949, n3425);
  not g6144 (n_2950, n3426);
  and g6145 (n3427, n_2949, n_2950);
  not g6146 (n_2951, n3427);
  and g6147 (n3428, n_2950, n_2951);
  not g6148 (n_2952, n3421);
  and g6149 (n3429, n_2952, n3428);
  and g6150 (n3430, n3423, n_2951);
  not g6151 (n_2953, n3429);
  not g6152 (n_2954, n3430);
  and g6153 (n3431, n_2953, n_2954);
  and g6154 (n3432, n1048, n1574);
  and g6155 (n3433, n891, n1919);
  and g6156 (n3434, \a[17] , \a[23] );
  and g6157 (n3435, n3165, n3434);
  not g6158 (n_2955, n3433);
  not g6159 (n_2956, n3435);
  and g6160 (n3436, n_2955, n_2956);
  not g6161 (n_2957, n3432);
  not g6162 (n_2958, n3436);
  and g6163 (n3437, n_2957, n_2958);
  not g6164 (n_2959, n3437);
  and g6165 (n3438, \a[23] , n_2959);
  and g6166 (n3439, \a[15] , n3438);
  and g6167 (n3440, \a[16] , \a[22] );
  and g6168 (n3441, \a[17] , \a[21] );
  not g6169 (n_2960, n3440);
  not g6170 (n_2961, n3441);
  and g6171 (n3442, n_2960, n_2961);
  and g6172 (n3443, n_2957, n_2959);
  not g6173 (n_2962, n3442);
  and g6174 (n3444, n_2962, n3443);
  not g6175 (n_2963, n3439);
  not g6176 (n_2964, n3444);
  and g6177 (n3445, n_2963, n_2964);
  not g6178 (n_2965, n3431);
  not g6179 (n_2966, n3445);
  and g6180 (n3446, n_2965, n_2966);
  not g6181 (n_2967, n3446);
  and g6182 (n3447, n_2965, n_2967);
  and g6183 (n3448, n_2966, n_2967);
  not g6184 (n_2968, n3447);
  not g6185 (n_2969, n3448);
  and g6186 (n3449, n_2968, n_2969);
  and g6187 (n3450, \a[9] , \a[29] );
  and g6188 (n3451, n380, n2865);
  and g6189 (n3452, \a[29] , \a[31] );
  and g6190 (n3453, n763, n3452);
  and g6191 (n3454, n432, n2617);
  not g6192 (n_2970, n3453);
  not g6193 (n_2971, n3454);
  and g6194 (n3455, n_2970, n_2971);
  not g6195 (n_2972, n3451);
  not g6196 (n_2973, n3455);
  and g6197 (n3456, n_2972, n_2973);
  not g6198 (n_2974, n3456);
  and g6199 (n3457, n3450, n_2974);
  and g6200 (n3458, n_2972, n_2974);
  and g6201 (n3459, \a[7] , \a[31] );
  and g6202 (n3460, \a[8] , \a[30] );
  not g6203 (n_2975, n3459);
  not g6204 (n_2976, n3460);
  and g6205 (n3461, n_2975, n_2976);
  not g6206 (n_2977, n3461);
  and g6207 (n3462, n3458, n_2977);
  not g6208 (n_2978, n3457);
  not g6209 (n_2979, n3462);
  and g6210 (n3463, n_2978, n_2979);
  not g6211 (n_2980, n3449);
  not g6212 (n_2981, n3463);
  and g6213 (n3464, n_2980, n_2981);
  not g6214 (n_2982, n3464);
  and g6215 (n3465, n_2980, n_2982);
  and g6216 (n3466, n_2981, n_2982);
  not g6217 (n_2983, n3465);
  not g6218 (n_2984, n3466);
  and g6219 (n3467, n_2983, n_2984);
  not g6220 (n_2985, n3467);
  and g6221 (n3468, n3418, n_2985);
  not g6222 (n_2986, n3418);
  and g6223 (n3469, n_2986, n3467);
  not g6224 (n_2987, n3408);
  not g6225 (n_2988, n3469);
  and g6226 (n3470, n_2987, n_2988);
  not g6227 (n_2989, n3468);
  and g6228 (n3471, n_2989, n3470);
  not g6229 (n_2990, n3471);
  and g6230 (n3472, n_2987, n_2990);
  and g6231 (n3473, n_2988, n_2990);
  and g6232 (n3474, n_2989, n3473);
  not g6233 (n_2991, n3472);
  not g6234 (n_2992, n3474);
  and g6235 (n3475, n_2991, n_2992);
  and g6236 (n3476, n_2805, n_2881);
  and g6237 (n3477, n3475, n3476);
  not g6238 (n_2993, n3475);
  not g6239 (n_2994, n3476);
  and g6240 (n3478, n_2993, n_2994);
  not g6241 (n_2995, n3477);
  not g6242 (n_2996, n3478);
  and g6243 (n3479, n_2995, n_2996);
  and g6244 (n3480, n_2904, n_2908);
  and g6245 (n3481, n_2771, n_2783);
  and g6246 (n3482, n_2857, n_2872);
  and g6247 (n3483, n3481, n3482);
  not g6248 (n_2997, n3481);
  not g6249 (n_2998, n3482);
  and g6250 (n3484, n_2997, n_2998);
  not g6251 (n_2999, n3483);
  not g6252 (n_3000, n3484);
  and g6253 (n3485, n_2999, n_3000);
  and g6254 (n3486, \a[1] , \a[37] );
  and g6255 (n3487, n1331, n3486);
  not g6256 (n_3001, n1331);
  not g6257 (n_3002, n3486);
  and g6258 (n3488, n_3001, n_3002);
  not g6259 (n_3003, n3487);
  not g6260 (n_3004, n3488);
  and g6261 (n3489, n_3003, n_3004);
  not g6262 (n_3005, n3489);
  and g6263 (n3490, n3286, n_3005);
  not g6264 (n_3006, n3286);
  and g6265 (n3491, n_3006, n3489);
  not g6266 (n_3007, n3490);
  not g6267 (n_3008, n3491);
  and g6268 (n3492, n_3007, n_3008);
  not g6269 (n_3009, n3341);
  and g6270 (n3493, n_3009, n3492);
  not g6271 (n_3010, n3492);
  and g6272 (n3494, n3341, n_3010);
  not g6273 (n_3011, n3493);
  not g6274 (n_3012, n3494);
  and g6275 (n3495, n_3011, n_3012);
  and g6276 (n3496, n3485, n3495);
  not g6277 (n_3013, n3485);
  not g6278 (n_3014, n3495);
  and g6279 (n3497, n_3013, n_3014);
  not g6280 (n_3015, n3496);
  not g6281 (n_3016, n3497);
  and g6282 (n3498, n_3015, n_3016);
  not g6283 (n_3017, n3498);
  and g6284 (n3499, n3480, n_3017);
  not g6285 (n_3018, n3480);
  and g6286 (n3500, n_3018, n3498);
  not g6287 (n_3019, n3499);
  not g6288 (n_3020, n3500);
  and g6289 (n3501, n_3019, n_3020);
  and g6290 (n3502, n_2887, n_2892);
  and g6291 (n3503, \a[27] , \a[34] );
  and g6292 (n3504, n649, n3503);
  and g6293 (n3505, n602, n2227);
  and g6294 (n3506, \a[12] , \a[34] );
  and g6295 (n3507, n2232, n3506);
  not g6296 (n_3021, n3505);
  not g6297 (n_3022, n3507);
  and g6298 (n3508, n_3021, n_3022);
  not g6299 (n_3023, n3504);
  not g6300 (n_3024, n3508);
  and g6301 (n3509, n_3023, n_3024);
  not g6302 (n_3025, n3509);
  and g6303 (n3510, \a[26] , n_3025);
  and g6304 (n3511, \a[12] , n3510);
  and g6305 (n3512, n_3023, n_3025);
  and g6306 (n3513, \a[4] , \a[34] );
  and g6307 (n3514, \a[11] , \a[27] );
  not g6308 (n_3026, n3513);
  not g6309 (n_3027, n3514);
  and g6310 (n3515, n_3026, n_3027);
  not g6311 (n_3028, n3515);
  and g6312 (n3516, n3512, n_3028);
  not g6313 (n_3029, n3511);
  not g6314 (n_3030, n3516);
  and g6315 (n3517, n_3029, n_3030);
  not g6316 (n_3031, n3502);
  not g6317 (n_3032, n3517);
  and g6318 (n3518, n_3031, n_3032);
  not g6319 (n_3033, n3518);
  and g6320 (n3519, n_3031, n_3033);
  and g6321 (n3520, n_3032, n_3033);
  not g6322 (n_3034, n3519);
  not g6323 (n_3035, n3520);
  and g6324 (n3521, n_3034, n_3035);
  and g6325 (n3522, n_2789, n_2793);
  and g6326 (n3523, n3521, n3522);
  not g6327 (n_3036, n3521);
  not g6328 (n_3037, n3522);
  and g6329 (n3524, n_3036, n_3037);
  not g6330 (n_3038, n3523);
  not g6331 (n_3039, n3524);
  and g6332 (n3525, n_3038, n_3039);
  and g6333 (n3526, n_2896, n_2900);
  and g6334 (n3527, \a[0] , \a[38] );
  and g6335 (n3528, \a[2] , \a[36] );
  not g6336 (n_3041, n3527);
  not g6337 (n_3042, n3528);
  and g6338 (n3529, n_3041, n_3042);
  and g6339 (n3530, \a[36] , \a[38] );
  and g6340 (n3531, n196, n3530);
  not g6341 (n_3043, n3529);
  not g6342 (n_3044, n3531);
  and g6343 (n3532, n_3043, n_3044);
  and g6344 (n3533, n3361, n3532);
  not g6345 (n_3045, n3533);
  and g6346 (n3534, n_3044, n_3045);
  and g6347 (n3535, n_3043, n3534);
  and g6348 (n3536, n3361, n_3045);
  not g6349 (n_3046, n3535);
  not g6350 (n_3047, n3536);
  and g6351 (n3537, n_3046, n_3047);
  not g6352 (n_3048, n3537);
  and g6353 (n3538, n3271, n_3048);
  not g6354 (n_3049, n3271);
  and g6355 (n3539, n_3049, n3537);
  not g6356 (n_3050, n3538);
  not g6357 (n_3051, n3539);
  and g6358 (n3540, n_3050, n_3051);
  and g6359 (n3541, \a[13] , \a[25] );
  and g6360 (n3542, \a[14] , \a[24] );
  not g6361 (n_3052, n3541);
  not g6362 (n_3053, n3542);
  and g6363 (n3543, n_3052, n_3053);
  and g6364 (n3544, n745, n1904);
  not g6365 (n_3054, n3544);
  not g6368 (n_3055, n3543);
  not g6370 (n_3056, n3547);
  and g6371 (n3548, \a[35] , n_3056);
  and g6372 (n3549, \a[3] , n3548);
  and g6373 (n3550, n_3054, n_3056);
  and g6374 (n3551, n_3055, n3550);
  not g6375 (n_3057, n3549);
  not g6376 (n_3058, n3551);
  and g6377 (n3552, n_3057, n_3058);
  not g6378 (n_3059, n3540);
  not g6379 (n_3060, n3552);
  and g6380 (n3553, n_3059, n_3060);
  and g6381 (n3554, n3540, n3552);
  not g6382 (n_3061, n3553);
  not g6383 (n_3062, n3554);
  and g6384 (n3555, n_3061, n_3062);
  not g6385 (n_3063, n3555);
  and g6386 (n3556, n3526, n_3063);
  not g6387 (n_3064, n3526);
  and g6388 (n3557, n_3064, n3555);
  not g6389 (n_3065, n3556);
  not g6390 (n_3066, n3557);
  and g6391 (n3558, n_3065, n_3066);
  and g6392 (n3559, n3525, n3558);
  not g6393 (n_3067, n3525);
  not g6394 (n_3068, n3558);
  and g6395 (n3560, n_3067, n_3068);
  not g6396 (n_3069, n3559);
  not g6397 (n_3070, n3560);
  and g6398 (n3561, n_3069, n_3070);
  and g6399 (n3562, n3501, n3561);
  not g6400 (n_3071, n3501);
  not g6401 (n_3072, n3561);
  and g6402 (n3563, n_3071, n_3072);
  not g6403 (n_3073, n3562);
  not g6404 (n_3074, n3563);
  and g6405 (n3564, n_3073, n_3074);
  not g6406 (n_3075, n3479);
  not g6407 (n_3076, n3564);
  and g6408 (n3565, n_3075, n_3076);
  and g6409 (n3566, n3479, n3564);
  not g6410 (n_3077, n3565);
  not g6411 (n_3078, n3566);
  and g6412 (n3567, n_3077, n_3078);
  not g6413 (n_3079, n3401);
  and g6414 (n3568, n_3079, n3567);
  not g6415 (n_3080, n3567);
  and g6416 (n3569, n3401, n_3080);
  not g6417 (n_3081, n3568);
  not g6418 (n_3082, n3569);
  and g6419 (n3570, n_3081, n_3082);
  and g6420 (n3571, n_2921, n_2924);
  not g6421 (n_3083, n3571);
  and g6422 (n3572, n_2920, n_3083);
  not g6423 (n_3084, n3570);
  and g6424 (n3573, n_3084, n3572);
  not g6425 (n_3085, n3572);
  and g6426 (n3574, n3570, n_3085);
  not g6427 (n_3086, n3573);
  not g6428 (n_3087, n3574);
  and g6429 (\asquared[39] , n_3086, n_3087);
  and g6430 (n3576, n_2996, n_3078);
  and g6431 (n3577, n_3020, n_3073);
  and g6432 (n3578, n_3066, n_3069);
  and g6433 (n3579, \a[0] , \a[39] );
  and g6434 (n3580, n3487, n3579);
  not g6435 (n_3089, n3580);
  and g6436 (n3581, n3487, n_3089);
  and g6437 (n3582, n_3003, n3579);
  not g6438 (n_3090, n3581);
  not g6439 (n_3091, n3582);
  and g6440 (n3583, n_3090, n_3091);
  and g6441 (n3584, \a[38] , n1203);
  not g6442 (n_3092, n3584);
  and g6443 (n3585, \a[20] , n_3092);
  and g6444 (n3586, \a[1] , n_3092);
  and g6445 (n3587, \a[38] , n3586);
  not g6446 (n_3093, n3585);
  not g6447 (n_3094, n3587);
  and g6448 (n3588, n_3093, n_3094);
  not g6449 (n_3095, n3583);
  not g6450 (n_3096, n3588);
  and g6451 (n3589, n_3095, n_3096);
  not g6452 (n_3097, n3589);
  and g6453 (n3590, n_3095, n_3097);
  and g6454 (n3591, n_3096, n_3097);
  not g6455 (n_3098, n3590);
  not g6456 (n_3099, n3591);
  and g6457 (n3592, n_3098, n_3099);
  and g6458 (n3593, n_3008, n_3011);
  and g6459 (n3594, n3592, n3593);
  not g6460 (n_3100, n3592);
  not g6461 (n_3101, n3593);
  and g6462 (n3595, n_3100, n_3101);
  not g6463 (n_3102, n3594);
  not g6464 (n_3103, n3595);
  and g6465 (n3596, n_3102, n_3103);
  and g6466 (n3597, n_2936, n_2940);
  not g6467 (n_3104, n3596);
  and g6468 (n3598, n_3104, n3597);
  not g6469 (n_3105, n3597);
  and g6470 (n3599, n3596, n_3105);
  not g6471 (n_3106, n3598);
  not g6472 (n_3107, n3599);
  and g6473 (n3600, n_3106, n_3107);
  and g6474 (n3601, n3534, n3550);
  not g6475 (n_3108, n3534);
  not g6476 (n_3109, n3550);
  and g6477 (n3602, n_3108, n_3109);
  not g6478 (n_3110, n3601);
  not g6479 (n_3111, n3602);
  and g6480 (n3603, n_3110, n_3111);
  not g6481 (n_3112, n3603);
  and g6482 (n3604, n3443, n_3112);
  not g6483 (n_3113, n3443);
  and g6484 (n3605, n_3113, n3603);
  not g6485 (n_3114, n3604);
  not g6486 (n_3115, n3605);
  and g6487 (n3606, n_3114, n_3115);
  and g6488 (n3607, n_2967, n_2982);
  and g6489 (n3608, n_3049, n_3048);
  not g6490 (n_3116, n3608);
  and g6491 (n3609, n_3061, n_3116);
  and g6492 (n3610, n3607, n3609);
  not g6493 (n_3117, n3607);
  not g6494 (n_3118, n3609);
  and g6495 (n3611, n_3117, n_3118);
  not g6496 (n_3119, n3610);
  not g6497 (n_3120, n3611);
  and g6498 (n3612, n_3119, n_3120);
  and g6499 (n3613, n3606, n3612);
  not g6500 (n_3121, n3606);
  not g6501 (n_3122, n3612);
  and g6502 (n3614, n_3121, n_3122);
  not g6503 (n_3123, n3613);
  not g6504 (n_3124, n3614);
  and g6505 (n3615, n_3123, n_3124);
  and g6506 (n3616, n3600, n3615);
  not g6507 (n_3125, n3600);
  not g6508 (n_3126, n3615);
  and g6509 (n3617, n_3125, n_3126);
  not g6510 (n_3127, n3616);
  not g6511 (n_3128, n3617);
  and g6512 (n3618, n_3127, n_3128);
  not g6513 (n_3129, n3578);
  and g6514 (n3619, n_3129, n3618);
  not g6515 (n_3130, n3618);
  and g6516 (n3620, n3578, n_3130);
  not g6517 (n_3131, n3619);
  not g6518 (n_3132, n3620);
  and g6519 (n3621, n_3131, n_3132);
  not g6520 (n_3133, n3621);
  and g6521 (n3622, n3577, n_3133);
  not g6522 (n_3134, n3577);
  and g6523 (n3623, n_3134, n3621);
  not g6524 (n_3135, n3622);
  not g6525 (n_3136, n3623);
  and g6526 (n3624, n_3135, n_3136);
  and g6527 (n3625, n_2930, n_2990);
  and g6528 (n3626, n3458, n3512);
  not g6529 (n_3137, n3458);
  not g6530 (n_3138, n3512);
  and g6531 (n3627, n_3137, n_3138);
  not g6532 (n_3139, n3626);
  not g6533 (n_3140, n3627);
  and g6534 (n3628, n_3139, n_3140);
  not g6535 (n_3141, n3628);
  and g6536 (n3629, n3428, n_3141);
  not g6537 (n_3142, n3428);
  and g6538 (n3630, n_3142, n3628);
  not g6539 (n_3143, n3629);
  not g6540 (n_3144, n3630);
  and g6541 (n3631, n_3143, n_3144);
  and g6542 (n3632, n_3033, n_3039);
  not g6543 (n_3145, n3631);
  and g6544 (n3633, n_3145, n3632);
  not g6545 (n_3146, n3632);
  and g6546 (n3634, n3631, n_3146);
  not g6547 (n_3147, n3633);
  not g6548 (n_3148, n3634);
  and g6549 (n3635, n_3147, n_3148);
  and g6550 (n3636, \a[4] , \a[35] );
  and g6551 (n3637, \a[12] , \a[27] );
  not g6552 (n_3149, n3636);
  not g6553 (n_3150, n3637);
  and g6554 (n3638, n_3149, n_3150);
  and g6555 (n3639, n3636, n3637);
  not g6556 (n_3151, n3639);
  not g6559 (n_3152, n3638);
  not g6561 (n_3153, n3642);
  and g6562 (n3643, n_3151, n_3153);
  and g6563 (n3644, n_3152, n3643);
  and g6564 (n3645, \a[22] , n_3153);
  and g6565 (n3646, \a[17] , n3645);
  not g6566 (n_3154, n3644);
  not g6567 (n_3155, n3646);
  and g6568 (n3647, n_3154, n_3155);
  and g6569 (n3648, \a[18] , \a[21] );
  not g6570 (n_3156, n1490);
  not g6571 (n_3157, n3648);
  and g6572 (n3649, n_3156, n_3157);
  and g6573 (n3650, n1149, n1494);
  not g6574 (n_3158, n3650);
  not g6577 (n_3159, n3649);
  not g6579 (n_3160, n3653);
  and g6580 (n3654, \a[31] , n_3160);
  and g6581 (n3655, \a[8] , n3654);
  and g6582 (n3656, n_3158, n_3160);
  and g6583 (n3657, n_3159, n3656);
  not g6584 (n_3161, n3655);
  not g6585 (n_3162, n3657);
  and g6586 (n3658, n_3161, n_3162);
  not g6587 (n_3163, n3647);
  not g6588 (n_3164, n3658);
  and g6589 (n3659, n_3163, n_3164);
  not g6590 (n_3165, n3659);
  and g6591 (n3660, n_3163, n_3165);
  and g6592 (n3661, n_3164, n_3165);
  not g6593 (n_3166, n3660);
  not g6594 (n_3167, n3661);
  and g6595 (n3662, n_3166, n_3167);
  and g6596 (n3663, \a[34] , n2768);
  and g6597 (n3664, \a[5] , \a[34] );
  and g6598 (n3665, n1976, n3664);
  and g6599 (n3666, n723, n2334);
  not g6600 (n_3168, n3665);
  not g6601 (n_3169, n3666);
  and g6602 (n3667, n_3168, n_3169);
  not g6603 (n_3170, n3663);
  not g6604 (n_3171, n3667);
  and g6605 (n3668, n_3170, n_3171);
  not g6606 (n_3172, n3668);
  and g6607 (n3669, n1976, n_3172);
  and g6608 (n3670, n_3170, n_3172);
  and g6609 (n3671, \a[10] , \a[29] );
  not g6610 (n_3173, n3664);
  not g6611 (n_3174, n3671);
  and g6612 (n3672, n_3173, n_3174);
  not g6613 (n_3175, n3672);
  and g6614 (n3673, n3670, n_3175);
  not g6615 (n_3176, n3669);
  not g6616 (n_3177, n3673);
  and g6617 (n3674, n_3176, n_3177);
  not g6618 (n_3178, n3662);
  not g6619 (n_3179, n3674);
  and g6620 (n3675, n_3178, n_3179);
  not g6621 (n_3180, n3675);
  and g6622 (n3676, n_3178, n_3180);
  and g6623 (n3677, n_3179, n_3180);
  not g6624 (n_3181, n3676);
  not g6625 (n_3182, n3677);
  and g6626 (n3678, n_3181, n_3182);
  not g6627 (n_3183, n3678);
  and g6628 (n3679, n3635, n_3183);
  not g6629 (n_3184, n3635);
  and g6630 (n3680, n_3184, n3678);
  not g6631 (n_3185, n3625);
  not g6632 (n_3186, n3680);
  and g6633 (n3681, n_3185, n_3186);
  not g6634 (n_3187, n3679);
  and g6635 (n3682, n_3187, n3681);
  not g6636 (n_3188, n3682);
  and g6637 (n3683, n_3185, n_3188);
  and g6638 (n3684, n_3186, n_3188);
  and g6639 (n3685, n_3187, n3684);
  not g6640 (n_3189, n3683);
  not g6641 (n_3190, n3685);
  and g6642 (n3686, n_3189, n_3190);
  and g6643 (n3687, \a[36] , \a[37] );
  and g6644 (n3688, n218, n3687);
  and g6645 (n3689, \a[13] , \a[37] );
  and g6646 (n3690, n1990, n3689);
  not g6647 (n_3191, n3688);
  not g6648 (n_3192, n3690);
  and g6649 (n3691, n_3191, n_3192);
  and g6650 (n3692, \a[3] , \a[36] );
  and g6651 (n3693, \a[13] , \a[26] );
  and g6652 (n3694, n3692, n3693);
  not g6653 (n_3193, n3691);
  not g6654 (n_3194, n3694);
  and g6655 (n3695, n_3193, n_3194);
  not g6656 (n_3195, n3695);
  and g6657 (n3696, n_3194, n_3195);
  not g6658 (n_3196, n3692);
  not g6659 (n_3197, n3693);
  and g6660 (n3697, n_3196, n_3197);
  not g6661 (n_3198, n3697);
  and g6662 (n3698, n3696, n_3198);
  and g6663 (n3699, \a[37] , n_3195);
  and g6664 (n3700, \a[2] , n3699);
  not g6665 (n_3199, n3698);
  not g6666 (n_3200, n3700);
  and g6667 (n3701, n_3199, n_3200);
  and g6668 (n3702, n891, n1666);
  and g6669 (n3703, n893, n1547);
  and g6670 (n3704, n895, n1904);
  not g6671 (n_3201, n3703);
  not g6672 (n_3202, n3704);
  and g6673 (n3705, n_3201, n_3202);
  not g6674 (n_3203, n3702);
  not g6675 (n_3204, n3705);
  and g6676 (n3706, n_3203, n_3204);
  not g6677 (n_3205, n3706);
  and g6678 (n3707, \a[25] , n_3205);
  and g6679 (n3708, \a[14] , n3707);
  and g6680 (n3709, n_3203, n_3205);
  and g6681 (n3710, \a[15] , \a[24] );
  and g6682 (n3711, \a[16] , \a[23] );
  not g6683 (n_3206, n3710);
  not g6684 (n_3207, n3711);
  and g6685 (n3712, n_3206, n_3207);
  not g6686 (n_3208, n3712);
  and g6687 (n3713, n3709, n_3208);
  not g6688 (n_3209, n3708);
  not g6689 (n_3210, n3713);
  and g6690 (n3714, n_3209, n_3210);
  not g6691 (n_3211, n3701);
  not g6692 (n_3212, n3714);
  and g6693 (n3715, n_3211, n_3212);
  not g6694 (n_3213, n3715);
  and g6695 (n3716, n_3211, n_3213);
  and g6696 (n3717, n_3212, n_3213);
  not g6697 (n_3214, n3716);
  not g6698 (n_3215, n3717);
  and g6699 (n3718, n_3214, n_3215);
  and g6700 (n3719, \a[6] , \a[33] );
  and g6701 (n3720, n763, n2488);
  and g6702 (n3721, n335, n3143);
  and g6703 (n3722, \a[9] , \a[30] );
  and g6704 (n3723, n3719, n3722);
  not g6705 (n_3216, n3721);
  not g6706 (n_3217, n3723);
  and g6707 (n3724, n_3216, n_3217);
  not g6708 (n_3218, n3720);
  not g6709 (n_3219, n3724);
  and g6710 (n3725, n_3218, n_3219);
  not g6711 (n_3220, n3725);
  and g6712 (n3726, n3719, n_3220);
  and g6713 (n3727, n_3218, n_3220);
  and g6714 (n3728, \a[7] , \a[32] );
  not g6715 (n_3221, n3722);
  not g6716 (n_3222, n3728);
  and g6717 (n3729, n_3221, n_3222);
  not g6718 (n_3223, n3729);
  and g6719 (n3730, n3727, n_3223);
  not g6720 (n_3224, n3726);
  not g6721 (n_3225, n3730);
  and g6722 (n3731, n_3224, n_3225);
  not g6723 (n_3226, n3718);
  not g6724 (n_3227, n3731);
  and g6725 (n3732, n_3226, n_3227);
  not g6726 (n_3228, n3732);
  and g6727 (n3733, n_3226, n_3228);
  and g6728 (n3734, n_3227, n_3228);
  not g6729 (n_3229, n3733);
  not g6730 (n_3230, n3734);
  and g6731 (n3735, n_3229, n_3230);
  and g6732 (n3736, n_3000, n_3015);
  and g6733 (n3737, n3735, n3736);
  not g6734 (n_3231, n3735);
  not g6735 (n_3232, n3736);
  and g6736 (n3738, n_3231, n_3232);
  not g6737 (n_3233, n3737);
  not g6738 (n_3234, n3738);
  and g6739 (n3739, n_3233, n_3234);
  and g6740 (n3740, n_2944, n_2989);
  not g6741 (n_3235, n3740);
  and g6742 (n3741, n3739, n_3235);
  not g6743 (n_3236, n3739);
  and g6744 (n3742, n_3236, n3740);
  not g6745 (n_3237, n3741);
  not g6746 (n_3238, n3742);
  and g6747 (n3743, n_3237, n_3238);
  and g6748 (n3744, n3686, n3743);
  not g6749 (n_3239, n3686);
  not g6750 (n_3240, n3743);
  and g6751 (n3745, n_3239, n_3240);
  not g6752 (n_3241, n3744);
  not g6753 (n_3242, n3745);
  and g6754 (n3746, n_3241, n_3242);
  not g6755 (n_3243, n3746);
  and g6756 (n3747, n3624, n_3243);
  not g6757 (n_3244, n3624);
  and g6758 (n3748, n_3244, n3746);
  not g6759 (n_3245, n3747);
  not g6760 (n_3246, n3748);
  and g6761 (n3749, n_3245, n_3246);
  not g6762 (n_3247, n3576);
  and g6763 (n3750, n_3247, n3749);
  not g6764 (n_3248, n3749);
  and g6765 (n3751, n3576, n_3248);
  not g6766 (n_3249, n3750);
  not g6767 (n_3250, n3751);
  and g6768 (n3752, n_3249, n_3250);
  and g6769 (n3753, n_3082, n_3085);
  not g6770 (n_3251, n3753);
  and g6771 (n3754, n_3081, n_3251);
  not g6772 (n_3252, n3752);
  and g6773 (n3755, n_3252, n3754);
  not g6774 (n_3253, n3754);
  and g6775 (n3756, n3752, n_3253);
  not g6776 (n_3254, n3755);
  not g6777 (n_3255, n3756);
  and g6778 (\asquared[40] , n_3254, n_3255);
  and g6779 (n3758, n_3250, n_3253);
  not g6780 (n_3256, n3758);
  and g6781 (n3759, n_3249, n_3256);
  and g6782 (n3760, n_3136, n_3245);
  and g6783 (n3761, n_3239, n3743);
  not g6784 (n_3257, n3761);
  and g6785 (n3762, n_3188, n_3257);
  and g6786 (n3763, n_3234, n_3237);
  and g6787 (n3764, n_3148, n_3187);
  and g6788 (n3765, n3670, n3696);
  not g6789 (n_3258, n3670);
  not g6790 (n_3259, n3696);
  and g6791 (n3766, n_3258, n_3259);
  not g6792 (n_3260, n3765);
  not g6793 (n_3261, n3766);
  and g6794 (n3767, n_3260, n_3261);
  not g6795 (n_3262, n3767);
  and g6796 (n3768, n3643, n_3262);
  not g6797 (n_3263, n3643);
  and g6798 (n3769, n_3263, n3767);
  not g6799 (n_3264, n3768);
  not g6800 (n_3265, n3769);
  and g6801 (n3770, n_3264, n_3265);
  and g6802 (n3771, n_3165, n_3180);
  and g6803 (n3772, n_3213, n_3228);
  and g6804 (n3773, n3771, n3772);
  not g6805 (n_3266, n3771);
  not g6806 (n_3267, n3772);
  and g6807 (n3774, n_3266, n_3267);
  not g6808 (n_3268, n3773);
  not g6809 (n_3269, n3774);
  and g6810 (n3775, n_3268, n_3269);
  and g6811 (n3776, n3770, n3775);
  not g6812 (n_3270, n3770);
  not g6813 (n_3271, n3775);
  and g6814 (n3777, n_3270, n_3271);
  not g6815 (n_3272, n3776);
  not g6816 (n_3273, n3777);
  and g6817 (n3778, n_3272, n_3273);
  not g6818 (n_3274, n3764);
  and g6819 (n3779, n_3274, n3778);
  not g6820 (n_3275, n3778);
  and g6821 (n3780, n3764, n_3275);
  not g6822 (n_3276, n3779);
  not g6823 (n_3277, n3780);
  and g6824 (n3781, n_3276, n_3277);
  not g6825 (n_3278, n3763);
  and g6826 (n3782, n_3278, n3781);
  not g6827 (n_3279, n3781);
  and g6828 (n3783, n3763, n_3279);
  not g6829 (n_3280, n3782);
  not g6830 (n_3281, n3783);
  and g6831 (n3784, n_3280, n_3281);
  not g6832 (n_3282, n3762);
  and g6833 (n3785, n_3282, n3784);
  not g6834 (n_3283, n3785);
  and g6835 (n3786, n3784, n_3283);
  and g6836 (n3787, n_3282, n_3283);
  not g6837 (n_3284, n3786);
  not g6838 (n_3285, n3787);
  and g6839 (n3788, n_3284, n_3285);
  and g6840 (n3789, n3709, n3727);
  not g6841 (n_3286, n3709);
  not g6842 (n_3287, n3727);
  and g6843 (n3790, n_3286, n_3287);
  not g6844 (n_3288, n3789);
  not g6845 (n_3289, n3790);
  and g6846 (n3791, n_3288, n_3289);
  and g6847 (n3792, n_3089, n_3097);
  not g6848 (n_3290, n3791);
  and g6849 (n3793, n_3290, n3792);
  not g6850 (n_3291, n3792);
  and g6851 (n3794, n3791, n_3291);
  not g6852 (n_3292, n3793);
  not g6853 (n_3293, n3794);
  and g6854 (n3795, n_3292, n_3293);
  and g6855 (n3796, n_3103, n_3107);
  not g6856 (n_3294, n3795);
  and g6857 (n3797, n_3294, n3796);
  not g6858 (n_3295, n3796);
  and g6859 (n3798, n3795, n_3295);
  not g6860 (n_3296, n3797);
  not g6861 (n_3297, n3798);
  and g6862 (n3799, n_3296, n_3297);
  and g6863 (n3800, \a[0] , \a[40] );
  and g6864 (n3801, \a[2] , \a[38] );
  not g6865 (n_3299, n3800);
  not g6866 (n_3300, n3801);
  and g6867 (n3802, n_3299, n_3300);
  and g6868 (n3803, \a[38] , \a[40] );
  and g6869 (n3804, n196, n3803);
  not g6870 (n_3301, n3802);
  not g6871 (n_3302, n3804);
  and g6872 (n3805, n_3301, n_3302);
  and g6873 (n3806, n1469, n3805);
  not g6874 (n_3303, n3806);
  and g6875 (n3807, n_3302, n_3303);
  and g6876 (n3808, n_3301, n3807);
  and g6877 (n3809, n1469, n_3303);
  not g6878 (n_3304, n3808);
  not g6879 (n_3305, n3809);
  and g6880 (n3810, n_3304, n_3305);
  and g6881 (n3811, \a[7] , \a[33] );
  and g6882 (n3812, \a[31] , \a[32] );
  and g6883 (n3813, n432, n3812);
  and g6884 (n3814, n763, n2598);
  and g6885 (n3815, n380, n3143);
  not g6886 (n_3306, n3814);
  not g6887 (n_3307, n3815);
  and g6888 (n3816, n_3306, n_3307);
  not g6889 (n_3308, n3813);
  not g6890 (n_3309, n3816);
  and g6891 (n3817, n_3308, n_3309);
  not g6892 (n_3310, n3817);
  and g6893 (n3818, n3811, n_3310);
  and g6894 (n3819, n_3308, n_3310);
  and g6895 (n3820, \a[8] , \a[32] );
  not g6896 (n_3311, n3091);
  not g6897 (n_3312, n3820);
  and g6898 (n3821, n_3311, n_3312);
  not g6899 (n_3313, n3821);
  and g6900 (n3822, n3819, n_3313);
  not g6901 (n_3314, n3818);
  not g6902 (n_3315, n3822);
  and g6903 (n3823, n_3314, n_3315);
  not g6904 (n_3316, n3810);
  not g6905 (n_3317, n3823);
  and g6906 (n3824, n_3316, n_3317);
  not g6907 (n_3318, n3824);
  and g6908 (n3825, n_3316, n_3318);
  and g6909 (n3826, n_3317, n_3318);
  not g6910 (n_3319, n3825);
  not g6911 (n_3320, n3826);
  and g6912 (n3827, n_3319, n_3320);
  and g6913 (n3828, \a[35] , \a[36] );
  and g6914 (n3829, n226, n3828);
  and g6915 (n3830, \a[12] , \a[36] );
  and g6916 (n3831, n2452, n3830);
  not g6917 (n_3321, n3829);
  not g6918 (n_3322, n3831);
  and g6919 (n3832, n_3321, n_3322);
  and g6920 (n3833, \a[5] , \a[35] );
  and g6921 (n3834, \a[12] , \a[28] );
  and g6922 (n3835, n3833, n3834);
  not g6923 (n_3323, n3832);
  not g6924 (n_3324, n3835);
  and g6925 (n3836, n_3323, n_3324);
  not g6926 (n_3325, n3836);
  and g6927 (n3837, \a[36] , n_3325);
  and g6928 (n3838, \a[4] , n3837);
  and g6929 (n3839, n_3324, n_3325);
  not g6930 (n_3326, n3833);
  not g6931 (n_3327, n3834);
  and g6932 (n3840, n_3326, n_3327);
  not g6933 (n_3328, n3840);
  and g6934 (n3841, n3839, n_3328);
  not g6935 (n_3329, n3838);
  not g6936 (n_3330, n3841);
  and g6937 (n3842, n_3329, n_3330);
  not g6938 (n_3331, n3827);
  not g6939 (n_3332, n3842);
  and g6940 (n3843, n_3331, n_3332);
  not g6941 (n_3333, n3843);
  and g6942 (n3844, n_3331, n_3333);
  and g6943 (n3845, n_3332, n_3333);
  not g6944 (n_3334, n3844);
  not g6945 (n_3335, n3845);
  and g6946 (n3846, n_3334, n_3335);
  not g6947 (n_3336, n3799);
  and g6948 (n3847, n_3336, n3846);
  not g6949 (n_3337, n3846);
  and g6950 (n3848, n3799, n_3337);
  not g6951 (n_3338, n3847);
  not g6952 (n_3339, n3848);
  and g6953 (n3849, n_3338, n_3339);
  and g6954 (n3850, n_3127, n_3131);
  not g6955 (n_3340, n3850);
  and g6956 (n3851, n3849, n_3340);
  not g6957 (n_3341, n3849);
  and g6958 (n3852, n_3341, n3850);
  not g6959 (n_3342, n3851);
  not g6960 (n_3343, n3852);
  and g6961 (n3853, n_3342, n_3343);
  and g6962 (n3854, \a[13] , \a[27] );
  and g6963 (n3855, \a[14] , \a[26] );
  not g6964 (n_3344, n3854);
  not g6965 (n_3345, n3855);
  and g6966 (n3856, n_3344, n_3345);
  and g6967 (n3857, n745, n2227);
  not g6968 (n_3346, n3857);
  not g6971 (n_3347, n3856);
  not g6973 (n_3348, n3860);
  and g6974 (n3861, n_3346, n_3348);
  and g6975 (n3862, n_3347, n3861);
  and g6976 (n3863, \a[37] , n_3348);
  and g6977 (n3864, \a[3] , n3863);
  not g6978 (n_3349, n3862);
  not g6979 (n_3350, n3864);
  and g6980 (n3865, n_3349, n_3350);
  and g6981 (n3866, n1048, n1666);
  and g6982 (n3867, n993, n1547);
  and g6983 (n3868, n891, n1904);
  not g6984 (n_3351, n3867);
  not g6985 (n_3352, n3868);
  and g6986 (n3869, n_3351, n_3352);
  not g6987 (n_3353, n3866);
  not g6988 (n_3354, n3869);
  and g6989 (n3870, n_3353, n_3354);
  not g6990 (n_3355, n3870);
  and g6991 (n3871, \a[25] , n_3355);
  and g6992 (n3872, \a[15] , n3871);
  and g6993 (n3873, n_3353, n_3355);
  and g6994 (n3874, \a[16] , \a[24] );
  not g6995 (n_3356, n3434);
  not g6996 (n_3357, n3874);
  and g6997 (n3875, n_3356, n_3357);
  not g6998 (n_3358, n3875);
  and g6999 (n3876, n3873, n_3358);
  not g7000 (n_3359, n3872);
  not g7001 (n_3360, n3876);
  and g7002 (n3877, n_3359, n_3360);
  not g7003 (n_3361, n3865);
  not g7004 (n_3362, n3877);
  and g7005 (n3878, n_3361, n_3362);
  not g7006 (n_3363, n3878);
  and g7007 (n3879, n_3361, n_3363);
  and g7008 (n3880, n_3362, n_3363);
  not g7009 (n_3364, n3879);
  not g7010 (n_3365, n3880);
  and g7011 (n3881, n_3364, n_3365);
  and g7012 (n3882, \a[6] , \a[34] );
  and g7013 (n3883, \a[10] , \a[30] );
  and g7014 (n3884, n3882, n3883);
  and g7015 (n3885, n723, n2617);
  and g7016 (n3886, \a[11] , \a[34] );
  and g7017 (n3887, n2928, n3886);
  not g7018 (n_3366, n3885);
  not g7019 (n_3367, n3887);
  and g7020 (n3888, n_3366, n_3367);
  not g7021 (n_3368, n3884);
  not g7022 (n_3369, n3888);
  and g7023 (n3889, n_3368, n_3369);
  not g7024 (n_3370, n3889);
  and g7025 (n3890, \a[29] , n_3370);
  and g7026 (n3891, \a[11] , n3890);
  and g7027 (n3892, n_3368, n_3370);
  not g7028 (n_3371, n3882);
  not g7029 (n_3372, n3883);
  and g7030 (n3893, n_3371, n_3372);
  not g7031 (n_3373, n3893);
  and g7032 (n3894, n3892, n_3373);
  not g7033 (n_3374, n3891);
  not g7034 (n_3375, n3894);
  and g7035 (n3895, n_3374, n_3375);
  not g7036 (n_3376, n3881);
  not g7037 (n_3377, n3895);
  and g7038 (n3896, n_3376, n_3377);
  not g7039 (n_3378, n3896);
  and g7040 (n3897, n_3376, n_3378);
  and g7041 (n3898, n_3377, n_3378);
  not g7042 (n_3379, n3897);
  not g7043 (n_3380, n3898);
  and g7044 (n3899, n_3379, n_3380);
  and g7045 (n3900, n_3120, n_3123);
  not g7046 (n_3381, n3899);
  not g7047 (n_3382, n3900);
  and g7048 (n3901, n_3381, n_3382);
  and g7049 (n3902, n3899, n3900);
  not g7050 (n_3383, n3901);
  not g7051 (n_3384, n3902);
  and g7052 (n3903, n_3383, n_3384);
  and g7053 (n3904, n_3140, n_3144);
  and g7054 (n3905, n_3111, n_3115);
  and g7055 (n3906, n3904, n3905);
  not g7056 (n_3385, n3904);
  not g7057 (n_3386, n3905);
  and g7058 (n3907, n_3385, n_3386);
  not g7059 (n_3387, n3906);
  not g7060 (n_3388, n3907);
  and g7061 (n3908, n_3387, n_3388);
  and g7062 (n3909, \a[1] , \a[39] );
  and g7063 (n3910, n1492, n3909);
  not g7064 (n_3389, n1492);
  not g7065 (n_3390, n3909);
  and g7066 (n3911, n_3389, n_3390);
  not g7067 (n_3391, n3910);
  not g7068 (n_3392, n3911);
  and g7069 (n3912, n_3391, n_3392);
  and g7070 (n3913, n3584, n3912);
  not g7071 (n_3393, n3912);
  and g7072 (n3914, n_3092, n_3393);
  not g7073 (n_3394, n3913);
  not g7074 (n_3395, n3914);
  and g7075 (n3915, n_3394, n_3395);
  not g7076 (n_3396, n3656);
  and g7077 (n3916, n_3396, n3915);
  not g7078 (n_3397, n3915);
  and g7079 (n3917, n3656, n_3397);
  not g7080 (n_3398, n3916);
  not g7081 (n_3399, n3917);
  and g7082 (n3918, n_3398, n_3399);
  and g7083 (n3919, n3908, n3918);
  not g7084 (n_3400, n3908);
  not g7085 (n_3401, n3918);
  and g7086 (n3920, n_3400, n_3401);
  not g7087 (n_3402, n3919);
  not g7088 (n_3403, n3920);
  and g7089 (n3921, n_3402, n_3403);
  and g7090 (n3922, n3903, n3921);
  not g7091 (n_3404, n3903);
  not g7092 (n_3405, n3921);
  and g7093 (n3923, n_3404, n_3405);
  not g7094 (n_3406, n3922);
  not g7095 (n_3407, n3923);
  and g7096 (n3924, n_3406, n_3407);
  and g7097 (n3925, n3853, n3924);
  not g7098 (n_3408, n3853);
  not g7099 (n_3409, n3924);
  and g7100 (n3926, n_3408, n_3409);
  not g7101 (n_3410, n3925);
  not g7102 (n_3411, n3926);
  and g7103 (n3927, n_3410, n_3411);
  not g7104 (n_3412, n3788);
  and g7105 (n3928, n_3412, n3927);
  not g7106 (n_3413, n3927);
  and g7107 (n3929, n_3285, n_3413);
  and g7108 (n3930, n_3284, n3929);
  not g7109 (n_3414, n3928);
  not g7110 (n_3415, n3930);
  and g7111 (n3931, n_3414, n_3415);
  not g7112 (n_3416, n3760);
  and g7113 (n3932, n_3416, n3931);
  not g7114 (n_3417, n3931);
  and g7115 (n3933, n3760, n_3417);
  not g7116 (n_3418, n3932);
  not g7117 (n_3419, n3933);
  and g7118 (n3934, n_3418, n_3419);
  not g7119 (n_3420, n3934);
  and g7120 (n3935, n3759, n_3420);
  not g7121 (n_3421, n3759);
  and g7122 (n3936, n_3421, n_3419);
  and g7123 (n3937, n_3418, n3936);
  not g7124 (n_3422, n3935);
  not g7125 (n_3423, n3937);
  and g7126 (\asquared[41] , n_3422, n_3423);
  and g7127 (n3939, n_3283, n_3414);
  and g7128 (n3940, n_3383, n_3406);
  and g7129 (n3941, n_3297, n_3339);
  and g7130 (n3942, n3807, n3873);
  not g7131 (n_3424, n3807);
  not g7132 (n_3425, n3873);
  and g7133 (n3943, n_3424, n_3425);
  not g7134 (n_3426, n3942);
  not g7135 (n_3427, n3943);
  and g7136 (n3944, n_3426, n_3427);
  not g7137 (n_3428, n3944);
  and g7138 (n3945, n3861, n_3428);
  not g7139 (n_3429, n3861);
  and g7140 (n3946, n_3429, n3944);
  not g7141 (n_3430, n3945);
  not g7142 (n_3431, n3946);
  and g7143 (n3947, n_3430, n_3431);
  and g7144 (n3948, n_3318, n_3333);
  not g7145 (n_3432, n3947);
  and g7146 (n3949, n_3432, n3948);
  not g7147 (n_3433, n3948);
  and g7148 (n3950, n3947, n_3433);
  not g7149 (n_3434, n3949);
  not g7150 (n_3435, n3950);
  and g7151 (n3951, n_3434, n_3435);
  and g7152 (n3952, \a[40] , n1296);
  and g7153 (n3953, \a[1] , \a[40] );
  not g7154 (n_3436, \a[21] );
  not g7155 (n_3437, n3953);
  and g7156 (n3954, n_3436, n_3437);
  not g7157 (n_3438, n3952);
  not g7158 (n_3439, n3954);
  and g7159 (n3955, n_3438, n_3439);
  not g7160 (n_3440, n3955);
  and g7161 (n3956, n3819, n_3440);
  not g7162 (n_3441, n3819);
  and g7163 (n3957, n_3441, n3955);
  not g7164 (n_3442, n3956);
  not g7165 (n_3443, n3957);
  and g7166 (n3958, n_3442, n_3443);
  not g7167 (n_3444, n3892);
  and g7168 (n3959, n_3444, n3958);
  not g7169 (n_3445, n3958);
  and g7170 (n3960, n3892, n_3445);
  not g7171 (n_3446, n3959);
  not g7172 (n_3447, n3960);
  and g7173 (n3961, n_3446, n_3447);
  and g7174 (n3962, n3951, n3961);
  not g7175 (n_3448, n3951);
  not g7176 (n_3449, n3961);
  and g7177 (n3963, n_3448, n_3449);
  not g7178 (n_3450, n3962);
  not g7179 (n_3451, n3963);
  and g7180 (n3964, n_3450, n_3451);
  not g7181 (n_3452, n3941);
  and g7182 (n3965, n_3452, n3964);
  not g7183 (n_3453, n3964);
  and g7184 (n3966, n3941, n_3453);
  not g7185 (n_3454, n3965);
  not g7186 (n_3455, n3966);
  and g7187 (n3967, n_3454, n_3455);
  not g7188 (n_3456, n3967);
  and g7189 (n3968, n3940, n_3456);
  not g7190 (n_3457, n3940);
  and g7191 (n3969, n_3457, n3967);
  not g7192 (n_3458, n3968);
  not g7193 (n_3459, n3969);
  and g7194 (n3970, n_3458, n_3459);
  and g7195 (n3971, n_3342, n_3410);
  not g7196 (n_3460, n3970);
  and g7197 (n3972, n_3460, n3971);
  not g7198 (n_3461, n3971);
  and g7199 (n3973, n3970, n_3461);
  not g7200 (n_3462, n3972);
  not g7201 (n_3463, n3973);
  and g7202 (n3974, n_3462, n_3463);
  and g7203 (n3975, n_3289, n_3293);
  and g7204 (n3976, n_3261, n_3265);
  and g7205 (n3977, n3975, n3976);
  not g7206 (n_3464, n3975);
  not g7207 (n_3465, n3976);
  and g7208 (n3978, n_3464, n_3465);
  not g7209 (n_3466, n3977);
  not g7210 (n_3467, n3978);
  and g7211 (n3979, n_3466, n_3467);
  and g7212 (n3980, n_3363, n_3378);
  not g7213 (n_3468, n3979);
  and g7214 (n3981, n_3468, n3980);
  not g7215 (n_3469, n3980);
  and g7216 (n3982, n3979, n_3469);
  not g7217 (n_3470, n3981);
  not g7218 (n_3471, n3982);
  and g7219 (n3983, n_3470, n_3471);
  and g7220 (n3984, \a[39] , \a[41] );
  and g7221 (n3985, n196, n3984);
  and g7222 (n3986, \a[0] , \a[41] );
  and g7223 (n3987, \a[2] , \a[39] );
  not g7224 (n_3473, n3986);
  not g7225 (n_3474, n3987);
  and g7226 (n3988, n_3473, n_3474);
  not g7227 (n_3475, n3985);
  not g7228 (n_3476, n3988);
  and g7229 (n3989, n_3475, n_3476);
  and g7230 (n3990, n3910, n3989);
  not g7231 (n_3477, n3989);
  and g7232 (n3991, n_3391, n_3477);
  not g7233 (n_3478, n3990);
  not g7234 (n_3479, n3991);
  and g7235 (n3992, n_3478, n_3479);
  not g7236 (n_3480, n3839);
  and g7237 (n3993, n_3480, n3992);
  not g7238 (n_3481, n3992);
  and g7239 (n3994, n3839, n_3481);
  not g7240 (n_3482, n3993);
  not g7241 (n_3483, n3994);
  and g7242 (n3995, n_3482, n_3483);
  and g7243 (n3996, \a[13] , \a[28] );
  and g7244 (n3997, \a[15] , \a[26] );
  not g7245 (n_3484, n3996);
  not g7246 (n_3485, n3997);
  and g7247 (n3998, n_3484, n_3485);
  and g7248 (n3999, n821, n2800);
  not g7249 (n_3486, n3999);
  not g7252 (n_3487, n3998);
  not g7254 (n_3488, n4002);
  and g7255 (n4003, \a[38] , n_3488);
  and g7256 (n4004, \a[3] , n4003);
  and g7257 (n4005, n_3486, n_3488);
  and g7258 (n4006, n_3487, n4005);
  not g7259 (n_3489, n4004);
  not g7260 (n_3490, n4006);
  and g7261 (n4007, n_3489, n_3490);
  not g7262 (n_3491, n4007);
  and g7263 (n4008, n3995, n_3491);
  not g7264 (n_3492, n4008);
  and g7265 (n4009, n3995, n_3492);
  and g7266 (n4010, n_3491, n_3492);
  not g7267 (n_3493, n4009);
  not g7268 (n_3494, n4010);
  and g7269 (n4011, n_3493, n_3494);
  and g7270 (n4012, n_3269, n_3272);
  not g7271 (n_3495, n4011);
  not g7272 (n_3496, n4012);
  and g7273 (n4013, n_3495, n_3496);
  not g7274 (n_3497, n4013);
  and g7275 (n4014, n_3495, n_3497);
  and g7276 (n4015, n_3496, n_3497);
  not g7277 (n_3498, n4014);
  not g7278 (n_3499, n4015);
  and g7279 (n4016, n_3498, n_3499);
  not g7280 (n_3500, n3983);
  and g7281 (n4017, n_3500, n4016);
  not g7282 (n_3501, n4016);
  and g7283 (n4018, n3983, n_3501);
  not g7284 (n_3502, n4017);
  not g7285 (n_3503, n4018);
  and g7286 (n4019, n_3502, n_3503);
  and g7287 (n4020, n_3276, n_3280);
  and g7288 (n4021, \a[6] , \a[35] );
  and g7289 (n4022, \a[11] , \a[30] );
  not g7290 (n_3504, n4021);
  not g7291 (n_3505, n4022);
  and g7292 (n4023, n_3504, n_3505);
  and g7293 (n4024, \a[30] , \a[35] );
  and g7294 (n4025, n815, n4024);
  and g7295 (n4026, n332, n3828);
  and g7296 (n4027, \a[30] , \a[36] );
  and g7297 (n4028, n502, n4027);
  not g7298 (n_3506, n4026);
  not g7299 (n_3507, n4028);
  and g7300 (n4029, n_3506, n_3507);
  not g7301 (n_3508, n4025);
  not g7302 (n_3509, n4029);
  and g7303 (n4030, n_3508, n_3509);
  not g7304 (n_3510, n4030);
  and g7305 (n4031, n_3508, n_3510);
  not g7306 (n_3511, n4023);
  and g7307 (n4032, n_3511, n4031);
  and g7308 (n4033, \a[36] , n_3510);
  and g7309 (n4034, \a[5] , n4033);
  not g7310 (n_3512, n4032);
  not g7311 (n_3513, n4034);
  and g7312 (n4035, n_3512, n_3513);
  and g7313 (n4036, \a[19] , \a[22] );
  not g7314 (n_3514, n1494);
  not g7315 (n_3515, n4036);
  and g7316 (n4037, n_3514, n_3515);
  and g7317 (n4038, n1494, n4036);
  not g7318 (n_3516, n4038);
  not g7321 (n_3517, n4037);
  not g7323 (n_3518, n4041);
  and g7324 (n4042, \a[33] , n_3518);
  and g7325 (n4043, \a[8] , n4042);
  and g7326 (n4044, n_3516, n_3518);
  and g7327 (n4045, n_3517, n4044);
  not g7328 (n_3519, n4043);
  not g7329 (n_3520, n4045);
  and g7330 (n4046, n_3519, n_3520);
  not g7331 (n_3521, n4035);
  not g7332 (n_3522, n4046);
  and g7333 (n4047, n_3521, n_3522);
  not g7334 (n_3523, n4047);
  and g7335 (n4048, n_3521, n_3523);
  and g7336 (n4049, n_3522, n_3523);
  not g7337 (n_3524, n4048);
  not g7338 (n_3525, n4049);
  and g7339 (n4050, n_3524, n_3525);
  and g7340 (n4051, n_3394, n_3398);
  and g7341 (n4052, n4050, n4051);
  not g7342 (n_3526, n4050);
  not g7343 (n_3527, n4051);
  and g7344 (n4053, n_3526, n_3527);
  not g7345 (n_3528, n4052);
  not g7346 (n_3529, n4053);
  and g7347 (n4054, n_3528, n_3529);
  and g7348 (n4055, n_3388, n_3402);
  not g7349 (n_3530, n4054);
  and g7350 (n4056, n_3530, n4055);
  not g7351 (n_3531, n4055);
  and g7352 (n4057, n4054, n_3531);
  not g7353 (n_3532, n4056);
  not g7354 (n_3533, n4057);
  and g7355 (n4058, n_3532, n_3533);
  and g7356 (n4059, \a[27] , \a[37] );
  and g7357 (n4060, n890, n4059);
  and g7358 (n4061, n606, n2041);
  not g7359 (n_3534, n4060);
  not g7360 (n_3535, n4061);
  and g7361 (n4062, n_3534, n_3535);
  and g7362 (n4063, \a[4] , \a[37] );
  and g7363 (n4064, \a[12] , \a[29] );
  and g7364 (n4065, n4063, n4064);
  not g7365 (n_3536, n4062);
  not g7366 (n_3537, n4065);
  and g7367 (n4066, n_3536, n_3537);
  not g7368 (n_3538, n4066);
  and g7369 (n4067, n_3537, n_3538);
  not g7370 (n_3539, n4063);
  not g7371 (n_3540, n4064);
  and g7372 (n4068, n_3539, n_3540);
  not g7373 (n_3541, n4068);
  and g7374 (n4069, n4067, n_3541);
  and g7375 (n4070, \a[27] , n_3538);
  and g7376 (n4071, \a[14] , n4070);
  not g7377 (n_3542, n4069);
  not g7378 (n_3543, n4071);
  and g7379 (n4072, n_3542, n_3543);
  and g7380 (n4073, n1052, n1666);
  and g7381 (n4074, n1050, n1547);
  and g7382 (n4075, n1048, n1904);
  not g7383 (n_3544, n4074);
  not g7384 (n_3545, n4075);
  and g7385 (n4076, n_3544, n_3545);
  not g7386 (n_3546, n4073);
  not g7387 (n_3547, n4076);
  and g7388 (n4077, n_3546, n_3547);
  not g7389 (n_3548, n4077);
  and g7390 (n4078, \a[25] , n_3548);
  and g7391 (n4079, \a[16] , n4078);
  and g7392 (n4080, n_3546, n_3548);
  and g7393 (n4081, \a[17] , \a[24] );
  and g7394 (n4082, \a[18] , \a[23] );
  not g7395 (n_3549, n4081);
  not g7396 (n_3550, n4082);
  and g7397 (n4083, n_3549, n_3550);
  not g7398 (n_3551, n4083);
  and g7399 (n4084, n4080, n_3551);
  not g7400 (n_3552, n4079);
  not g7401 (n_3553, n4084);
  and g7402 (n4085, n_3552, n_3553);
  not g7403 (n_3554, n4072);
  not g7404 (n_3555, n4085);
  and g7405 (n4086, n_3554, n_3555);
  not g7406 (n_3556, n4086);
  and g7407 (n4087, n_3554, n_3556);
  and g7408 (n4088, n_3555, n_3556);
  not g7409 (n_3557, n4087);
  not g7410 (n_3558, n4088);
  and g7411 (n4089, n_3557, n_3558);
  and g7412 (n4090, \a[32] , \a[34] );
  and g7413 (n4091, n763, n4090);
  and g7414 (n4092, n484, n3812);
  and g7415 (n4093, \a[7] , \a[34] );
  and g7416 (n4094, n2352, n4093);
  not g7417 (n_3559, n4092);
  not g7418 (n_3560, n4094);
  and g7419 (n4095, n_3559, n_3560);
  not g7420 (n_3561, n4091);
  not g7421 (n_3562, n4095);
  and g7422 (n4096, n_3561, n_3562);
  not g7423 (n_3563, n4096);
  and g7424 (n4097, n2352, n_3563);
  and g7425 (n4098, n_3561, n_3563);
  and g7426 (n4099, \a[9] , \a[32] );
  not g7427 (n_3564, n4093);
  not g7428 (n_3565, n4099);
  and g7429 (n4100, n_3564, n_3565);
  not g7430 (n_3566, n4100);
  and g7431 (n4101, n4098, n_3566);
  not g7432 (n_3567, n4097);
  not g7433 (n_3568, n4101);
  and g7434 (n4102, n_3567, n_3568);
  not g7435 (n_3569, n4089);
  not g7436 (n_3570, n4102);
  and g7437 (n4103, n_3569, n_3570);
  not g7438 (n_3571, n4103);
  and g7439 (n4104, n_3569, n_3571);
  and g7440 (n4105, n_3570, n_3571);
  not g7441 (n_3572, n4104);
  not g7442 (n_3573, n4105);
  and g7443 (n4106, n_3572, n_3573);
  not g7444 (n_3574, n4058);
  and g7445 (n4107, n_3574, n4106);
  not g7446 (n_3575, n4106);
  and g7447 (n4108, n4058, n_3575);
  not g7448 (n_3576, n4107);
  not g7449 (n_3577, n4108);
  and g7450 (n4109, n_3576, n_3577);
  not g7451 (n_3578, n4020);
  and g7452 (n4110, n_3578, n4109);
  not g7453 (n_3579, n4110);
  and g7454 (n4111, n_3578, n_3579);
  and g7455 (n4112, n4109, n_3579);
  not g7456 (n_3580, n4111);
  not g7457 (n_3581, n4112);
  and g7458 (n4113, n_3580, n_3581);
  not g7459 (n_3582, n4113);
  and g7460 (n4114, n4019, n_3582);
  not g7461 (n_3583, n4019);
  and g7462 (n4115, n_3583, n_3581);
  and g7463 (n4116, n_3580, n4115);
  not g7464 (n_3584, n4114);
  not g7465 (n_3585, n4116);
  and g7466 (n4117, n_3584, n_3585);
  and g7467 (n4118, n3974, n4117);
  not g7468 (n_3586, n3974);
  not g7469 (n_3587, n4117);
  and g7470 (n4119, n_3586, n_3587);
  not g7471 (n_3588, n4118);
  not g7472 (n_3589, n4119);
  and g7473 (n4120, n_3588, n_3589);
  not g7474 (n_3590, n4120);
  and g7475 (n4121, n3939, n_3590);
  not g7476 (n_3591, n3939);
  and g7477 (n4122, n_3591, n4120);
  not g7478 (n_3592, n4121);
  not g7479 (n_3593, n4122);
  and g7480 (n4123, n_3592, n_3593);
  not g7481 (n_3594, n3936);
  and g7482 (n4124, n_3418, n_3594);
  not g7483 (n_3595, n4123);
  and g7484 (n4125, n_3595, n4124);
  not g7485 (n_3596, n4124);
  and g7486 (n4126, n4123, n_3596);
  not g7487 (n_3597, n4125);
  not g7488 (n_3598, n4126);
  and g7489 (\asquared[42] , n_3597, n_3598);
  and g7490 (n4128, n_3592, n_3596);
  not g7491 (n_3599, n4128);
  and g7492 (n4129, n_3593, n_3599);
  and g7493 (n4130, n_3463, n_3588);
  and g7494 (n4131, n_3454, n_3459);
  and g7495 (n4132, n_3467, n_3471);
  and g7496 (n4133, \a[7] , \a[35] );
  and g7497 (n4134, \a[11] , \a[31] );
  and g7498 (n4135, n4133, n4134);
  and g7499 (n4136, \a[31] , \a[36] );
  and g7500 (n4137, n815, n4136);
  and g7501 (n4138, n335, n3828);
  not g7502 (n_3600, n4137);
  not g7503 (n_3601, n4138);
  and g7504 (n4139, n_3600, n_3601);
  not g7505 (n_3602, n4135);
  not g7506 (n_3603, n4139);
  and g7507 (n4140, n_3602, n_3603);
  not g7508 (n_3604, n4140);
  and g7509 (n4141, \a[6] , n_3604);
  and g7510 (n4142, \a[36] , n4141);
  and g7511 (n4143, n_3602, n_3604);
  not g7512 (n_3605, n4133);
  not g7513 (n_3606, n4134);
  and g7514 (n4144, n_3605, n_3606);
  not g7515 (n_3607, n4144);
  and g7516 (n4145, n4143, n_3607);
  not g7517 (n_3608, n4142);
  not g7518 (n_3609, n4145);
  and g7519 (n4146, n_3608, n_3609);
  not g7520 (n_3610, n4146);
  and g7521 (n4147, n4098, n_3610);
  not g7522 (n_3611, n4098);
  and g7523 (n4148, n_3611, n4146);
  not g7524 (n_3612, n4147);
  not g7525 (n_3613, n4148);
  and g7526 (n4149, n_3612, n_3613);
  and g7527 (n4150, \a[33] , \a[34] );
  and g7528 (n4151, n432, n4150);
  and g7529 (n4152, n378, n4090);
  and g7530 (n4153, n484, n3143);
  not g7531 (n_3614, n4152);
  not g7532 (n_3615, n4153);
  and g7533 (n4154, n_3614, n_3615);
  not g7534 (n_3616, n4151);
  not g7535 (n_3617, n4154);
  and g7536 (n4155, n_3616, n_3617);
  not g7537 (n_3618, n4155);
  and g7538 (n4156, n3264, n_3618);
  and g7539 (n4157, n_3616, n_3618);
  and g7540 (n4158, \a[8] , \a[34] );
  and g7541 (n4159, \a[9] , \a[33] );
  not g7542 (n_3619, n4158);
  not g7543 (n_3620, n4159);
  and g7544 (n4160, n_3619, n_3620);
  not g7545 (n_3621, n4160);
  and g7546 (n4161, n4157, n_3621);
  not g7547 (n_3622, n4156);
  not g7548 (n_3623, n4161);
  and g7549 (n4162, n_3622, n_3623);
  not g7550 (n_3624, n4149);
  not g7551 (n_3625, n4162);
  and g7552 (n4163, n_3624, n_3625);
  and g7553 (n4164, n4149, n4162);
  not g7554 (n_3626, n4163);
  not g7555 (n_3627, n4164);
  and g7556 (n4165, n_3626, n_3627);
  not g7557 (n_3628, n4165);
  and g7558 (n4166, n4132, n_3628);
  not g7559 (n_3629, n4132);
  and g7560 (n4167, n_3629, n4165);
  not g7561 (n_3630, n4166);
  not g7562 (n_3631, n4167);
  and g7563 (n4168, n_3630, n_3631);
  and g7564 (n4169, \a[16] , \a[40] );
  and g7565 (n4170, n1990, n4169);
  and g7566 (n4171, \a[39] , \a[40] );
  and g7567 (n4172, n218, n4171);
  not g7568 (n_3632, n4170);
  not g7569 (n_3633, n4172);
  and g7570 (n4173, n_3632, n_3633);
  and g7571 (n4174, \a[3] , \a[39] );
  and g7572 (n4175, \a[16] , \a[26] );
  and g7573 (n4176, n4174, n4175);
  not g7574 (n_3634, n4173);
  not g7575 (n_3635, n4176);
  and g7576 (n4177, n_3634, n_3635);
  not g7577 (n_3636, n4177);
  and g7578 (n4178, n_3635, n_3636);
  not g7579 (n_3637, n4174);
  not g7580 (n_3638, n4175);
  and g7581 (n4179, n_3637, n_3638);
  not g7582 (n_3639, n4179);
  and g7583 (n4180, n4178, n_3639);
  and g7584 (n4181, \a[40] , n_3636);
  and g7585 (n4182, \a[2] , n4181);
  not g7586 (n_3640, n4180);
  not g7587 (n_3641, n4182);
  and g7588 (n4183, n_3640, n_3641);
  and g7589 (n4184, n1149, n1666);
  and g7590 (n4185, n1547, n3134);
  and g7591 (n4186, n1052, n1904);
  not g7592 (n_3642, n4185);
  not g7593 (n_3643, n4186);
  and g7594 (n4187, n_3642, n_3643);
  not g7595 (n_3644, n4184);
  not g7596 (n_3645, n4187);
  and g7597 (n4188, n_3644, n_3645);
  not g7598 (n_3646, n4188);
  and g7599 (n4189, \a[25] , n_3646);
  and g7600 (n4190, \a[17] , n4189);
  and g7601 (n4191, \a[18] , \a[24] );
  and g7602 (n4192, \a[19] , \a[23] );
  not g7603 (n_3647, n4191);
  not g7604 (n_3648, n4192);
  and g7605 (n4193, n_3647, n_3648);
  and g7606 (n4194, n_3644, n_3646);
  not g7607 (n_3649, n4193);
  and g7608 (n4195, n_3649, n4194);
  not g7609 (n_3650, n4190);
  not g7610 (n_3651, n4195);
  and g7611 (n4196, n_3650, n_3651);
  not g7612 (n_3652, n4183);
  not g7613 (n_3653, n4196);
  and g7614 (n4197, n_3652, n_3653);
  not g7615 (n_3654, n4197);
  and g7616 (n4198, n_3652, n_3654);
  and g7617 (n4199, n_3653, n_3654);
  not g7618 (n_3655, n4198);
  not g7619 (n_3656, n4199);
  and g7620 (n4200, n_3655, n_3656);
  and g7621 (n4201, \a[14] , \a[38] );
  and g7622 (n4202, n2452, n4201);
  and g7623 (n4203, n895, n2331);
  and g7624 (n4204, \a[15] , \a[38] );
  and g7625 (n4205, n2341, n4204);
  not g7626 (n_3657, n4203);
  not g7627 (n_3658, n4205);
  and g7628 (n4206, n_3657, n_3658);
  not g7629 (n_3659, n4202);
  not g7630 (n_3660, n4206);
  and g7631 (n4207, n_3659, n_3660);
  not g7632 (n_3661, n4207);
  and g7633 (n4208, \a[27] , n_3661);
  and g7634 (n4209, \a[15] , n4208);
  and g7635 (n4210, n_3659, n_3661);
  and g7636 (n4211, \a[4] , \a[38] );
  and g7637 (n4212, \a[14] , \a[28] );
  not g7638 (n_3662, n4211);
  not g7639 (n_3663, n4212);
  and g7640 (n4213, n_3662, n_3663);
  not g7641 (n_3664, n4213);
  and g7642 (n4214, n4210, n_3664);
  not g7643 (n_3665, n4209);
  not g7644 (n_3666, n4214);
  and g7645 (n4215, n_3665, n_3666);
  not g7646 (n_3667, n4200);
  not g7647 (n_3668, n4215);
  and g7648 (n4216, n_3667, n_3668);
  not g7649 (n_3669, n4216);
  and g7650 (n4217, n_3667, n_3669);
  and g7651 (n4218, n_3668, n_3669);
  not g7652 (n_3670, n4217);
  not g7653 (n_3671, n4218);
  and g7654 (n4219, n_3670, n_3671);
  not g7655 (n_3672, n4219);
  and g7656 (n4220, n4168, n_3672);
  not g7657 (n_3673, n4168);
  and g7658 (n4221, n_3673, n4219);
  not g7659 (n_3674, n4131);
  not g7660 (n_3675, n4221);
  and g7661 (n4222, n_3674, n_3675);
  not g7662 (n_3676, n4220);
  and g7663 (n4223, n_3676, n4222);
  not g7664 (n_3677, n4223);
  and g7665 (n4224, n_3674, n_3677);
  and g7666 (n4225, n_3675, n_3677);
  and g7667 (n4226, n_3676, n4225);
  not g7668 (n_3678, n4224);
  not g7669 (n_3679, n4226);
  and g7670 (n4227, n_3678, n_3679);
  and g7671 (n4228, \a[0] , \a[42] );
  and g7672 (n4229, n3952, n4228);
  not g7673 (n_3681, n4229);
  and g7674 (n4230, n3952, n_3681);
  and g7675 (n4231, n_3438, n4228);
  not g7676 (n_3682, n4230);
  not g7677 (n_3683, n4231);
  and g7678 (n4232, n_3682, n_3683);
  and g7679 (n4233, \a[1] , \a[41] );
  and g7680 (n4234, n1693, n4233);
  not g7681 (n_3684, n4234);
  and g7682 (n4235, n4233, n_3684);
  and g7683 (n4236, n1693, n_3684);
  not g7684 (n_3685, n4235);
  not g7685 (n_3686, n4236);
  and g7686 (n4237, n_3685, n_3686);
  not g7687 (n_3687, n4232);
  not g7688 (n_3688, n4237);
  and g7689 (n4238, n_3687, n_3688);
  not g7690 (n_3689, n4238);
  and g7691 (n4239, n_3687, n_3689);
  and g7692 (n4240, n_3688, n_3689);
  not g7693 (n_3690, n4239);
  not g7694 (n_3691, n4240);
  and g7695 (n4241, n_3690, n_3691);
  and g7696 (n4242, \a[5] , \a[37] );
  and g7697 (n4243, \a[12] , \a[30] );
  and g7698 (n4244, n4242, n4243);
  and g7699 (n4245, n748, n2617);
  and g7700 (n4246, n2772, n3689);
  not g7701 (n_3692, n4245);
  not g7702 (n_3693, n4246);
  and g7703 (n4247, n_3692, n_3693);
  not g7704 (n_3694, n4244);
  not g7705 (n_3695, n4247);
  and g7706 (n4248, n_3694, n_3695);
  not g7707 (n_3696, n4248);
  and g7708 (n4249, \a[29] , n_3696);
  and g7709 (n4250, \a[13] , n4249);
  and g7710 (n4251, n_3694, n_3696);
  not g7711 (n_3697, n4242);
  not g7712 (n_3698, n4243);
  and g7713 (n4252, n_3697, n_3698);
  not g7714 (n_3699, n4252);
  and g7715 (n4253, n4251, n_3699);
  not g7716 (n_3700, n4250);
  not g7717 (n_3701, n4253);
  and g7718 (n4254, n_3700, n_3701);
  not g7719 (n_3702, n4241);
  not g7720 (n_3703, n4254);
  and g7721 (n4255, n_3702, n_3703);
  not g7722 (n_3704, n4255);
  and g7723 (n4256, n_3702, n_3704);
  and g7724 (n4257, n_3703, n_3704);
  not g7725 (n_3705, n4256);
  not g7726 (n_3706, n4257);
  and g7727 (n4258, n_3705, n_3706);
  and g7728 (n4259, n_3443, n_3446);
  and g7729 (n4260, n4258, n4259);
  not g7730 (n_3707, n4258);
  not g7731 (n_3708, n4259);
  and g7732 (n4261, n_3707, n_3708);
  not g7733 (n_3709, n4260);
  not g7734 (n_3710, n4261);
  and g7735 (n4262, n_3709, n_3710);
  and g7736 (n4263, n_3435, n_3450);
  not g7737 (n_3711, n4262);
  and g7738 (n4264, n_3711, n4263);
  not g7739 (n_3712, n4263);
  and g7740 (n4265, n4262, n_3712);
  not g7741 (n_3713, n4264);
  not g7742 (n_3714, n4265);
  and g7743 (n4266, n_3713, n_3714);
  and g7744 (n4267, n4044, n4067);
  not g7745 (n_3715, n4044);
  not g7746 (n_3716, n4067);
  and g7747 (n4268, n_3715, n_3716);
  not g7748 (n_3717, n4267);
  not g7749 (n_3718, n4268);
  and g7750 (n4269, n_3717, n_3718);
  not g7751 (n_3719, n4269);
  and g7752 (n4270, n4031, n_3719);
  not g7753 (n_3720, n4031);
  and g7754 (n4271, n_3720, n4269);
  not g7755 (n_3721, n4270);
  not g7756 (n_3722, n4271);
  and g7757 (n4272, n_3721, n_3722);
  and g7758 (n4273, n_3523, n_3529);
  not g7759 (n_3723, n4272);
  and g7760 (n4274, n_3723, n4273);
  not g7761 (n_3724, n4273);
  and g7762 (n4275, n4272, n_3724);
  not g7763 (n_3725, n4274);
  not g7764 (n_3726, n4275);
  and g7765 (n4276, n_3725, n_3726);
  and g7766 (n4277, n4005, n4080);
  not g7767 (n_3727, n4005);
  not g7768 (n_3728, n4080);
  and g7769 (n4278, n_3727, n_3728);
  not g7770 (n_3729, n4277);
  not g7771 (n_3730, n4278);
  and g7772 (n4279, n_3729, n_3730);
  and g7773 (n4280, n_3475, n_3478);
  not g7774 (n_3731, n4279);
  and g7775 (n4281, n_3731, n4280);
  not g7776 (n_3732, n4280);
  and g7777 (n4282, n4279, n_3732);
  not g7778 (n_3733, n4281);
  not g7779 (n_3734, n4282);
  and g7780 (n4283, n_3733, n_3734);
  and g7781 (n4284, n4276, n4283);
  not g7782 (n_3735, n4276);
  not g7783 (n_3736, n4283);
  and g7784 (n4285, n_3735, n_3736);
  not g7785 (n_3737, n4284);
  not g7786 (n_3738, n4285);
  and g7787 (n4286, n_3737, n_3738);
  and g7788 (n4287, n4266, n4286);
  not g7789 (n_3739, n4266);
  not g7790 (n_3740, n4286);
  and g7791 (n4288, n_3739, n_3740);
  not g7792 (n_3741, n4287);
  not g7793 (n_3742, n4288);
  and g7794 (n4289, n_3741, n_3742);
  and g7795 (n4290, n4227, n4289);
  not g7796 (n_3743, n4227);
  not g7797 (n_3744, n4289);
  and g7798 (n4291, n_3743, n_3744);
  not g7799 (n_3745, n4290);
  not g7800 (n_3746, n4291);
  and g7801 (n4292, n_3745, n_3746);
  and g7802 (n4293, n_3579, n_3584);
  and g7803 (n4294, n_3497, n_3503);
  and g7804 (n4295, n_3427, n_3431);
  and g7805 (n4296, n_3482, n_3492);
  and g7806 (n4297, n4295, n4296);
  not g7807 (n_3747, n4295);
  not g7808 (n_3748, n4296);
  and g7809 (n4298, n_3747, n_3748);
  not g7810 (n_3749, n4297);
  not g7811 (n_3750, n4298);
  and g7812 (n4299, n_3749, n_3750);
  and g7813 (n4300, n_3556, n_3571);
  not g7814 (n_3751, n4299);
  and g7815 (n4301, n_3751, n4300);
  not g7816 (n_3752, n4300);
  and g7817 (n4302, n4299, n_3752);
  not g7818 (n_3753, n4301);
  not g7819 (n_3754, n4302);
  and g7820 (n4303, n_3753, n_3754);
  and g7821 (n4304, n_3533, n_3577);
  not g7822 (n_3755, n4304);
  and g7823 (n4305, n4303, n_3755);
  not g7824 (n_3756, n4303);
  and g7825 (n4306, n_3756, n4304);
  not g7826 (n_3757, n4305);
  not g7827 (n_3758, n4306);
  and g7828 (n4307, n_3757, n_3758);
  not g7829 (n_3759, n4294);
  and g7830 (n4308, n_3759, n4307);
  not g7831 (n_3760, n4307);
  and g7832 (n4309, n4294, n_3760);
  not g7833 (n_3761, n4308);
  not g7834 (n_3762, n4309);
  and g7835 (n4310, n_3761, n_3762);
  not g7836 (n_3763, n4293);
  and g7837 (n4311, n_3763, n4310);
  not g7838 (n_3764, n4310);
  and g7839 (n4312, n4293, n_3764);
  not g7840 (n_3765, n4311);
  not g7841 (n_3766, n4312);
  and g7842 (n4313, n_3765, n_3766);
  not g7843 (n_3767, n4292);
  and g7844 (n4314, n_3767, n4313);
  not g7845 (n_3768, n4314);
  and g7846 (n4315, n4313, n_3768);
  and g7847 (n4316, n_3767, n_3768);
  not g7848 (n_3769, n4315);
  not g7849 (n_3770, n4316);
  and g7850 (n4317, n_3769, n_3770);
  not g7851 (n_3771, n4130);
  not g7852 (n_3772, n4317);
  and g7853 (n4318, n_3771, n_3772);
  and g7854 (n4319, n4130, n4317);
  not g7855 (n_3773, n4318);
  not g7856 (n_3774, n4319);
  and g7857 (n4320, n_3773, n_3774);
  not g7858 (n_3775, n4129);
  and g7859 (n4321, n_3775, n4320);
  not g7860 (n_3776, n4320);
  and g7861 (n4322, n4129, n_3776);
  not g7862 (n_3777, n4321);
  not g7863 (n_3778, n4322);
  and g7864 (\asquared[43] , n_3777, n_3778);
  and g7865 (n4324, n_3765, n_3768);
  and g7866 (n4325, n_3743, n4289);
  not g7867 (n_3779, n4325);
  and g7868 (n4326, n_3677, n_3779);
  and g7869 (n4327, n_3714, n_3741);
  and g7870 (n4328, n_3631, n_3676);
  and g7871 (n4329, n_3654, n_3669);
  and g7872 (n4330, n_3611, n_3610);
  not g7873 (n_3780, n4330);
  and g7874 (n4331, n_3626, n_3780);
  and g7875 (n4332, \a[42] , n1405);
  and g7876 (n4333, \a[1] , \a[42] );
  not g7877 (n_3781, \a[22] );
  not g7878 (n_3782, n4333);
  and g7879 (n4334, n_3781, n_3782);
  not g7880 (n_3783, n4332);
  not g7881 (n_3784, n4334);
  and g7882 (n4335, n_3783, n_3784);
  and g7883 (n4336, n4234, n4335);
  not g7884 (n_3785, n4335);
  and g7885 (n4337, n_3684, n_3785);
  not g7886 (n_3786, n4336);
  not g7887 (n_3787, n4337);
  and g7888 (n4338, n_3786, n_3787);
  not g7889 (n_3788, n4157);
  and g7890 (n4339, n_3788, n4338);
  not g7891 (n_3789, n4338);
  and g7892 (n4340, n4157, n_3789);
  not g7893 (n_3790, n4339);
  not g7894 (n_3791, n4340);
  and g7895 (n4341, n_3790, n_3791);
  not g7896 (n_3792, n4331);
  and g7897 (n4342, n_3792, n4341);
  not g7898 (n_3793, n4342);
  and g7899 (n4343, n_3792, n_3793);
  and g7900 (n4344, n4341, n_3793);
  not g7901 (n_3794, n4343);
  not g7902 (n_3795, n4344);
  and g7903 (n4345, n_3794, n_3795);
  not g7904 (n_3796, n4329);
  not g7905 (n_3797, n4345);
  and g7906 (n4346, n_3796, n_3797);
  and g7907 (n4347, n4329, n_3795);
  and g7908 (n4348, n_3794, n4347);
  not g7909 (n_3798, n4346);
  not g7910 (n_3799, n4348);
  and g7911 (n4349, n_3798, n_3799);
  not g7912 (n_3800, n4328);
  and g7913 (n4350, n_3800, n4349);
  not g7914 (n_3801, n4349);
  and g7915 (n4351, n4328, n_3801);
  not g7916 (n_3802, n4350);
  not g7917 (n_3803, n4351);
  and g7918 (n4352, n_3802, n_3803);
  not g7919 (n_3804, n4327);
  and g7920 (n4353, n_3804, n4352);
  not g7921 (n_3805, n4352);
  and g7922 (n4354, n4327, n_3805);
  not g7923 (n_3806, n4353);
  not g7924 (n_3807, n4354);
  and g7925 (n4355, n_3806, n_3807);
  not g7926 (n_3808, n4326);
  and g7927 (n4356, n_3808, n4355);
  not g7928 (n_3809, n4356);
  and g7929 (n4357, n_3808, n_3809);
  and g7930 (n4358, n4355, n_3809);
  not g7931 (n_3810, n4357);
  not g7932 (n_3811, n4358);
  and g7933 (n4359, n_3810, n_3811);
  and g7934 (n4360, n_3757, n_3761);
  and g7935 (n4361, n_3750, n_3754);
  and g7936 (n4362, n209, n4171);
  and g7937 (n4363, \a[4] , \a[43] );
  and g7938 (n4364, n3579, n4363);
  not g7939 (n_3813, n4362);
  not g7940 (n_3814, n4364);
  and g7941 (n4365, n_3813, n_3814);
  and g7942 (n4366, \a[0] , \a[43] );
  and g7943 (n4367, \a[3] , \a[40] );
  and g7944 (n4368, n4366, n4367);
  not g7945 (n_3815, n4365);
  not g7946 (n_3816, n4368);
  and g7947 (n4369, n_3815, n_3816);
  not g7948 (n_3817, n4369);
  and g7949 (n4370, n_3816, n_3817);
  not g7950 (n_3818, n4366);
  not g7951 (n_3819, n4367);
  and g7952 (n4371, n_3818, n_3819);
  not g7953 (n_3820, n4371);
  and g7954 (n4372, n4370, n_3820);
  and g7955 (n4373, \a[39] , n_3817);
  and g7956 (n4374, \a[4] , n4373);
  not g7957 (n_3821, n4372);
  not g7958 (n_3822, n4374);
  and g7959 (n4375, n_3821, n_3822);
  and g7960 (n4376, n891, n2331);
  and g7961 (n4377, n893, n2041);
  and g7962 (n4378, n895, n2334);
  not g7963 (n_3823, n4377);
  not g7964 (n_3824, n4378);
  and g7965 (n4379, n_3823, n_3824);
  not g7966 (n_3825, n4376);
  not g7967 (n_3826, n4379);
  and g7968 (n4380, n_3825, n_3826);
  not g7969 (n_3827, n4380);
  and g7970 (n4381, \a[29] , n_3827);
  and g7971 (n4382, \a[14] , n4381);
  and g7972 (n4383, n_3825, n_3827);
  and g7973 (n4384, \a[15] , \a[28] );
  and g7974 (n4385, \a[16] , \a[27] );
  not g7975 (n_3828, n4384);
  not g7976 (n_3829, n4385);
  and g7977 (n4386, n_3828, n_3829);
  not g7978 (n_3830, n4386);
  and g7979 (n4387, n4383, n_3830);
  not g7980 (n_3831, n4382);
  not g7981 (n_3832, n4387);
  and g7982 (n4388, n_3831, n_3832);
  not g7983 (n_3833, n4375);
  not g7984 (n_3834, n4388);
  and g7985 (n4389, n_3833, n_3834);
  not g7986 (n_3835, n4389);
  and g7987 (n4390, n_3833, n_3835);
  and g7988 (n4391, n_3834, n_3835);
  not g7989 (n_3836, n4390);
  not g7990 (n_3837, n4391);
  and g7991 (n4392, n_3836, n_3837);
  and g7992 (n4393, n1149, n1904);
  and g7993 (n4394, n2301, n3134);
  and g7994 (n4395, n1052, n2463);
  not g7995 (n_3838, n4394);
  not g7996 (n_3839, n4395);
  and g7997 (n4396, n_3838, n_3839);
  not g7998 (n_3840, n4393);
  not g7999 (n_3841, n4396);
  and g8000 (n4397, n_3840, n_3841);
  not g8001 (n_3842, n4397);
  and g8002 (n4398, \a[26] , n_3842);
  and g8003 (n4399, \a[17] , n4398);
  and g8004 (n4400, \a[18] , \a[25] );
  not g8005 (n_3843, n1664);
  not g8006 (n_3844, n4400);
  and g8007 (n4401, n_3843, n_3844);
  and g8008 (n4402, n_3840, n_3842);
  not g8009 (n_3845, n4401);
  and g8010 (n4403, n_3845, n4402);
  not g8011 (n_3846, n4399);
  not g8012 (n_3847, n4403);
  and g8013 (n4404, n_3846, n_3847);
  not g8014 (n_3848, n4392);
  not g8015 (n_3849, n4404);
  and g8016 (n4405, n_3848, n_3849);
  not g8017 (n_3850, n4405);
  and g8018 (n4406, n_3848, n_3850);
  and g8019 (n4407, n_3849, n_3850);
  not g8020 (n_3851, n4406);
  not g8021 (n_3852, n4407);
  and g8022 (n4408, n_3851, n_3852);
  and g8023 (n4409, n378, n2972);
  and g8024 (n4410, n380, n3828);
  and g8025 (n4411, \a[10] , \a[36] );
  and g8026 (n4412, n3811, n4411);
  not g8027 (n_3853, n4410);
  not g8028 (n_3854, n4412);
  and g8029 (n4413, n_3853, n_3854);
  not g8030 (n_3855, n4409);
  not g8031 (n_3856, n4413);
  and g8032 (n4414, n_3855, n_3856);
  not g8033 (n_3857, n4414);
  and g8034 (n4415, n_3855, n_3857);
  and g8035 (n4416, \a[8] , \a[35] );
  and g8036 (n4417, \a[10] , \a[33] );
  not g8037 (n_3858, n4416);
  not g8038 (n_3859, n4417);
  and g8039 (n4418, n_3858, n_3859);
  not g8040 (n_3860, n4418);
  and g8041 (n4419, n4415, n_3860);
  and g8042 (n4420, \a[36] , n_3857);
  and g8043 (n4421, \a[7] , n4420);
  not g8044 (n_3861, n4419);
  not g8045 (n_3862, n4421);
  and g8046 (n4422, n_3861, n_3862);
  and g8047 (n4423, \a[20] , \a[23] );
  not g8048 (n_3863, n1574);
  not g8049 (n_3864, n4423);
  and g8050 (n4424, n_3863, n_3864);
  and g8051 (n4425, n1494, n1919);
  not g8052 (n_3865, n4425);
  not g8055 (n_3866, n4424);
  not g8057 (n_3867, n4428);
  and g8058 (n4429, \a[34] , n_3867);
  and g8059 (n4430, \a[9] , n4429);
  and g8060 (n4431, n_3865, n_3867);
  and g8061 (n4432, n_3866, n4431);
  not g8062 (n_3868, n4430);
  not g8063 (n_3869, n4432);
  and g8064 (n4433, n_3868, n_3869);
  not g8065 (n_3870, n4422);
  not g8066 (n_3871, n4433);
  and g8067 (n4434, n_3870, n_3871);
  not g8068 (n_3872, n4434);
  and g8069 (n4435, n_3870, n_3872);
  and g8070 (n4436, n_3871, n_3872);
  not g8071 (n_3873, n4435);
  not g8072 (n_3874, n4436);
  and g8073 (n4437, n_3873, n_3874);
  and g8074 (n4438, \a[5] , \a[38] );
  and g8075 (n4439, \a[13] , \a[30] );
  not g8076 (n_3875, n4438);
  not g8077 (n_3876, n4439);
  and g8078 (n4440, n_3875, n_3876);
  and g8079 (n4441, n4438, n4439);
  not g8080 (n_3877, n4441);
  not g8083 (n_3878, n4440);
  not g8085 (n_3879, n4444);
  and g8086 (n4445, \a[41] , n_3879);
  and g8087 (n4446, \a[2] , n4445);
  and g8088 (n4447, n_3877, n_3879);
  and g8089 (n4448, n_3878, n4447);
  not g8090 (n_3880, n4446);
  not g8091 (n_3881, n4448);
  and g8092 (n4449, n_3880, n_3881);
  not g8093 (n_3882, n4437);
  not g8094 (n_3883, n4449);
  and g8095 (n4450, n_3882, n_3883);
  not g8096 (n_3884, n4450);
  and g8097 (n4451, n_3882, n_3884);
  and g8098 (n4452, n_3883, n_3884);
  not g8099 (n_3885, n4451);
  not g8100 (n_3886, n4452);
  and g8101 (n4453, n_3885, n_3886);
  not g8102 (n_3887, n4408);
  and g8103 (n4454, n_3887, n4453);
  not g8104 (n_3888, n4453);
  and g8105 (n4455, n4408, n_3888);
  not g8106 (n_3889, n4454);
  not g8107 (n_3890, n4455);
  and g8108 (n4456, n_3889, n_3890);
  not g8109 (n_3891, n4361);
  not g8110 (n_3892, n4456);
  and g8111 (n4457, n_3891, n_3892);
  and g8112 (n4458, n4361, n4456);
  not g8113 (n_3893, n4457);
  not g8114 (n_3894, n4458);
  and g8115 (n4459, n_3893, n_3894);
  not g8116 (n_3895, n4360);
  and g8117 (n4460, n_3895, n4459);
  not g8118 (n_3896, n4459);
  and g8119 (n4461, n4360, n_3896);
  not g8120 (n_3897, n4460);
  not g8121 (n_3898, n4461);
  and g8122 (n4462, n_3897, n_3898);
  and g8123 (n4463, n_3704, n_3710);
  and g8124 (n4464, n4143, n4210);
  not g8125 (n_3899, n4143);
  not g8126 (n_3900, n4210);
  and g8127 (n4465, n_3899, n_3900);
  not g8128 (n_3901, n4464);
  not g8129 (n_3902, n4465);
  and g8130 (n4466, n_3901, n_3902);
  not g8131 (n_3903, n4466);
  and g8132 (n4467, n4194, n_3903);
  not g8133 (n_3904, n4194);
  and g8134 (n4468, n_3904, n4466);
  not g8135 (n_3905, n4467);
  not g8136 (n_3906, n4468);
  and g8137 (n4469, n_3905, n_3906);
  and g8138 (n4470, n4178, n4251);
  not g8139 (n_3907, n4178);
  not g8140 (n_3908, n4251);
  and g8141 (n4471, n_3907, n_3908);
  not g8142 (n_3909, n4470);
  not g8143 (n_3910, n4471);
  and g8144 (n4472, n_3909, n_3910);
  and g8145 (n4473, n_3681, n_3689);
  not g8146 (n_3911, n4472);
  and g8147 (n4474, n_3911, n4473);
  not g8148 (n_3912, n4473);
  and g8149 (n4475, n4472, n_3912);
  not g8150 (n_3913, n4474);
  not g8151 (n_3914, n4475);
  and g8152 (n4476, n_3913, n_3914);
  not g8153 (n_3915, n4469);
  not g8154 (n_3916, n4476);
  and g8155 (n4477, n_3915, n_3916);
  and g8156 (n4478, n4469, n4476);
  not g8157 (n_3917, n4477);
  not g8158 (n_3918, n4478);
  and g8159 (n4479, n_3917, n_3918);
  not g8160 (n_3919, n4463);
  and g8161 (n4480, n_3919, n4479);
  not g8162 (n_3920, n4479);
  and g8163 (n4481, n4463, n_3920);
  not g8164 (n_3921, n4480);
  not g8165 (n_3922, n4481);
  and g8166 (n4482, n_3921, n_3922);
  and g8167 (n4483, n_3718, n_3722);
  and g8168 (n4484, n602, n3812);
  and g8169 (n4485, \a[12] , \a[37] );
  and g8170 (n4486, n3336, n4485);
  not g8171 (n_3923, n4484);
  not g8172 (n_3924, n4486);
  and g8173 (n4487, n_3923, n_3924);
  and g8174 (n4488, \a[6] , \a[37] );
  and g8175 (n4489, \a[11] , \a[32] );
  and g8176 (n4490, n4488, n4489);
  not g8177 (n_3925, n4487);
  not g8178 (n_3926, n4490);
  and g8179 (n4491, n_3925, n_3926);
  not g8180 (n_3927, n4491);
  and g8181 (n4492, \a[31] , n_3927);
  and g8182 (n4493, \a[12] , n4492);
  and g8183 (n4494, n_3926, n_3927);
  not g8184 (n_3928, n4488);
  not g8185 (n_3929, n4489);
  and g8186 (n4495, n_3928, n_3929);
  not g8187 (n_3930, n4495);
  and g8188 (n4496, n4494, n_3930);
  not g8189 (n_3931, n4493);
  not g8190 (n_3932, n4496);
  and g8191 (n4497, n_3931, n_3932);
  not g8192 (n_3933, n4483);
  not g8193 (n_3934, n4497);
  and g8194 (n4498, n_3933, n_3934);
  not g8195 (n_3935, n4498);
  and g8196 (n4499, n_3933, n_3935);
  and g8197 (n4500, n_3934, n_3935);
  not g8198 (n_3936, n4499);
  not g8199 (n_3937, n4500);
  and g8200 (n4501, n_3936, n_3937);
  and g8201 (n4502, n_3730, n_3734);
  and g8202 (n4503, n4501, n4502);
  not g8203 (n_3938, n4501);
  not g8204 (n_3939, n4502);
  and g8205 (n4504, n_3938, n_3939);
  not g8206 (n_3940, n4503);
  not g8207 (n_3941, n4504);
  and g8208 (n4505, n_3940, n_3941);
  and g8209 (n4506, n_3726, n_3737);
  not g8210 (n_3942, n4506);
  and g8211 (n4507, n4505, n_3942);
  not g8212 (n_3943, n4505);
  and g8213 (n4508, n_3943, n4506);
  not g8214 (n_3944, n4507);
  not g8215 (n_3945, n4508);
  and g8216 (n4509, n_3944, n_3945);
  and g8217 (n4510, n4482, n4509);
  not g8218 (n_3946, n4482);
  not g8219 (n_3947, n4509);
  and g8220 (n4511, n_3946, n_3947);
  not g8221 (n_3948, n4510);
  not g8222 (n_3949, n4511);
  and g8223 (n4512, n_3948, n_3949);
  and g8224 (n4513, n4462, n4512);
  not g8225 (n_3950, n4462);
  not g8226 (n_3951, n4512);
  and g8227 (n4514, n_3950, n_3951);
  not g8228 (n_3952, n4513);
  not g8229 (n_3953, n4514);
  and g8230 (n4515, n_3952, n_3953);
  not g8231 (n_3954, n4359);
  and g8232 (n4516, n_3954, n4515);
  not g8233 (n_3955, n4515);
  and g8234 (n4517, n_3811, n_3955);
  and g8235 (n4518, n_3810, n4517);
  not g8236 (n_3956, n4516);
  not g8237 (n_3957, n4518);
  and g8238 (n4519, n_3956, n_3957);
  not g8239 (n_3958, n4324);
  and g8240 (n4520, n_3958, n4519);
  not g8241 (n_3959, n4519);
  and g8242 (n4521, n4324, n_3959);
  not g8243 (n_3960, n4520);
  not g8244 (n_3961, n4521);
  and g8245 (n4522, n_3960, n_3961);
  and g8246 (n4523, n_3775, n_3774);
  not g8247 (n_3962, n4523);
  and g8248 (n4524, n_3773, n_3962);
  not g8249 (n_3963, n4522);
  and g8250 (n4525, n_3963, n4524);
  not g8251 (n_3964, n4524);
  and g8252 (n4526, n4522, n_3964);
  not g8253 (n_3965, n4525);
  not g8254 (n_3966, n4526);
  and g8255 (\asquared[44] , n_3965, n_3966);
  and g8256 (n4528, n_3809, n_3956);
  and g8257 (n4529, n_3802, n_3806);
  and g8258 (n4530, n_3793, n_3798);
  and g8259 (n4531, \a[15] , \a[29] );
  and g8260 (n4532, \a[17] , \a[27] );
  not g8261 (n_3967, n4531);
  not g8262 (n_3968, n4532);
  and g8263 (n4533, n_3967, n_3968);
  and g8264 (n4534, n993, n2041);
  not g8265 (n_3969, n4534);
  not g8268 (n_3970, n4533);
  not g8270 (n_3971, n4537);
  and g8271 (n4538, n_3969, n_3971);
  and g8272 (n4539, n_3970, n4538);
  and g8273 (n4540, \a[41] , n_3971);
  and g8274 (n4541, \a[3] , n4540);
  not g8275 (n_3972, n4539);
  not g8276 (n_3973, n4541);
  and g8277 (n4542, n_3972, n_3973);
  and g8278 (n4543, \a[18] , \a[26] );
  and g8279 (n4544, n1490, n1904);
  and g8280 (n4545, n1331, n2301);
  and g8281 (n4546, n1149, n2463);
  not g8282 (n_3974, n4545);
  not g8283 (n_3975, n4546);
  and g8284 (n4547, n_3974, n_3975);
  not g8285 (n_3976, n4544);
  not g8286 (n_3977, n4547);
  and g8287 (n4548, n_3976, n_3977);
  not g8288 (n_3978, n4548);
  and g8289 (n4549, n4543, n_3978);
  and g8290 (n4550, \a[19] , \a[25] );
  and g8291 (n4551, \a[20] , \a[24] );
  not g8292 (n_3979, n4550);
  not g8293 (n_3980, n4551);
  and g8294 (n4552, n_3979, n_3980);
  and g8295 (n4553, n_3976, n_3978);
  not g8296 (n_3981, n4552);
  and g8297 (n4554, n_3981, n4553);
  not g8298 (n_3982, n4549);
  not g8299 (n_3983, n4554);
  and g8300 (n4555, n_3982, n_3983);
  not g8301 (n_3984, n4542);
  not g8302 (n_3985, n4555);
  and g8303 (n4556, n_3984, n_3985);
  not g8304 (n_3986, n4556);
  and g8305 (n4557, n_3984, n_3986);
  and g8306 (n4558, n_3985, n_3986);
  not g8307 (n_3987, n4557);
  not g8308 (n_3988, n4558);
  and g8309 (n4559, n_3987, n_3988);
  and g8310 (n4560, \a[6] , \a[38] );
  and g8311 (n4561, \a[11] , \a[37] );
  and g8312 (n4562, n3811, n4561);
  and g8313 (n4563, \a[33] , \a[38] );
  and g8314 (n4564, n815, n4563);
  and g8315 (n4565, \a[37] , \a[38] );
  and g8316 (n4566, n335, n4565);
  not g8317 (n_3989, n4564);
  not g8318 (n_3990, n4566);
  and g8319 (n4567, n_3989, n_3990);
  not g8320 (n_3991, n4562);
  not g8321 (n_3992, n4567);
  and g8322 (n4568, n_3991, n_3992);
  not g8323 (n_3993, n4568);
  and g8324 (n4569, n4560, n_3993);
  and g8325 (n4570, n_3991, n_3993);
  and g8326 (n4571, \a[7] , \a[37] );
  and g8327 (n4572, \a[11] , \a[33] );
  not g8328 (n_3994, n4571);
  not g8329 (n_3995, n4572);
  and g8330 (n4573, n_3994, n_3995);
  not g8331 (n_3996, n4573);
  and g8332 (n4574, n4570, n_3996);
  not g8333 (n_3997, n4569);
  not g8334 (n_3998, n4574);
  and g8335 (n4575, n_3997, n_3998);
  not g8336 (n_3999, n4559);
  not g8337 (n_4000, n4575);
  and g8338 (n4576, n_3999, n_4000);
  not g8339 (n_4001, n4576);
  and g8340 (n4577, n_3999, n_4001);
  and g8341 (n4578, n_4000, n_4001);
  not g8342 (n_4002, n4577);
  not g8343 (n_4003, n4578);
  and g8344 (n4579, n_4002, n_4003);
  and g8345 (n4580, n2452, n4169);
  and g8346 (n4581, n893, n3110);
  not g8347 (n_4004, n4580);
  not g8348 (n_4005, n4581);
  and g8349 (n4582, n_4004, n_4005);
  and g8350 (n4583, \a[4] , \a[40] );
  and g8351 (n4584, \a[14] , \a[30] );
  and g8352 (n4585, n4583, n4584);
  not g8353 (n_4006, n4582);
  not g8354 (n_4007, n4585);
  and g8355 (n4586, n_4006, n_4007);
  not g8356 (n_4008, n4586);
  and g8357 (n4587, n_4007, n_4008);
  not g8358 (n_4009, n4583);
  not g8359 (n_4010, n4584);
  and g8360 (n4588, n_4009, n_4010);
  not g8361 (n_4011, n4588);
  and g8362 (n4589, n4587, n_4011);
  and g8363 (n4590, \a[28] , n_4008);
  and g8364 (n4591, \a[16] , n4590);
  not g8365 (n_4012, n4589);
  not g8366 (n_4013, n4591);
  and g8367 (n4592, n_4012, n_4013);
  and g8368 (n4593, \a[8] , \a[36] );
  and g8369 (n4594, n484, n3319);
  and g8370 (n4595, \a[34] , \a[36] );
  and g8371 (n4596, n378, n4595);
  and g8372 (n4597, n432, n3828);
  not g8373 (n_4014, n4596);
  not g8374 (n_4015, n4597);
  and g8375 (n4598, n_4014, n_4015);
  not g8376 (n_4016, n4594);
  not g8377 (n_4017, n4598);
  and g8378 (n4599, n_4016, n_4017);
  not g8379 (n_4018, n4599);
  and g8380 (n4600, n4593, n_4018);
  and g8381 (n4601, n_4016, n_4018);
  and g8382 (n4602, \a[9] , \a[35] );
  and g8383 (n4603, \a[10] , \a[34] );
  not g8384 (n_4019, n4602);
  not g8385 (n_4020, n4603);
  and g8386 (n4604, n_4019, n_4020);
  not g8387 (n_4021, n4604);
  and g8388 (n4605, n4601, n_4021);
  not g8389 (n_4022, n4600);
  not g8390 (n_4023, n4605);
  and g8391 (n4606, n_4022, n_4023);
  not g8392 (n_4024, n4592);
  not g8393 (n_4025, n4606);
  and g8394 (n4607, n_4024, n_4025);
  not g8395 (n_4026, n4607);
  and g8396 (n4608, n_4024, n_4026);
  and g8397 (n4609, n_4025, n_4026);
  not g8398 (n_4027, n4608);
  not g8399 (n_4028, n4609);
  and g8400 (n4610, n_4027, n_4028);
  and g8401 (n4611, \a[12] , \a[32] );
  and g8402 (n4612, \a[13] , \a[31] );
  not g8403 (n_4029, n4611);
  not g8404 (n_4030, n4612);
  and g8405 (n4613, n_4029, n_4030);
  and g8406 (n4614, n748, n3812);
  not g8407 (n_4031, n4614);
  not g8410 (n_4032, n4613);
  not g8412 (n_4033, n4617);
  and g8413 (n4618, \a[39] , n_4033);
  and g8414 (n4619, \a[5] , n4618);
  and g8415 (n4620, n_4031, n_4033);
  and g8416 (n4621, n_4032, n4620);
  not g8417 (n_4034, n4619);
  not g8418 (n_4035, n4621);
  and g8419 (n4622, n_4034, n_4035);
  not g8420 (n_4036, n4610);
  not g8421 (n_4037, n4622);
  and g8422 (n4623, n_4036, n_4037);
  not g8423 (n_4038, n4623);
  and g8424 (n4624, n_4036, n_4038);
  and g8425 (n4625, n_4037, n_4038);
  not g8426 (n_4039, n4624);
  not g8427 (n_4040, n4625);
  and g8428 (n4626, n_4039, n_4040);
  and g8429 (n4627, n4579, n4626);
  not g8430 (n_4041, n4579);
  not g8431 (n_4042, n4626);
  and g8432 (n4628, n_4041, n_4042);
  not g8433 (n_4043, n4627);
  not g8434 (n_4044, n4628);
  and g8435 (n4629, n_4043, n_4044);
  not g8436 (n_4045, n4530);
  and g8437 (n4630, n_4045, n4629);
  not g8438 (n_4046, n4629);
  and g8439 (n4631, n4530, n_4046);
  not g8440 (n_4047, n4630);
  not g8441 (n_4048, n4631);
  and g8442 (n4632, n_4047, n_4048);
  not g8443 (n_4049, n4632);
  and g8444 (n4633, n4529, n_4049);
  not g8445 (n_4050, n4529);
  and g8446 (n4634, n_4050, n4632);
  not g8447 (n_4051, n4633);
  not g8448 (n_4052, n4634);
  and g8449 (n4635, n_4051, n_4052);
  and g8450 (n4636, n4383, n4494);
  not g8451 (n_4053, n4383);
  not g8452 (n_4054, n4494);
  and g8453 (n4637, n_4053, n_4054);
  not g8454 (n_4055, n4636);
  not g8455 (n_4056, n4637);
  and g8456 (n4638, n_4055, n_4056);
  and g8457 (n4639, \a[42] , \a[44] );
  and g8458 (n4640, n196, n4639);
  and g8459 (n4641, \a[0] , \a[44] );
  and g8460 (n4642, \a[2] , \a[42] );
  not g8461 (n_4058, n4641);
  not g8462 (n_4059, n4642);
  and g8463 (n4643, n_4058, n_4059);
  not g8464 (n_4060, n4640);
  not g8465 (n_4061, n4643);
  and g8466 (n4644, n_4060, n_4061);
  and g8467 (n4645, n4332, n4644);
  not g8468 (n_4062, n4645);
  and g8469 (n4646, n4332, n_4062);
  and g8470 (n4647, n_4060, n_4062);
  and g8471 (n4648, n_4061, n4647);
  not g8472 (n_4063, n4646);
  not g8473 (n_4064, n4648);
  and g8474 (n4649, n_4063, n_4064);
  not g8475 (n_4065, n4649);
  and g8476 (n4650, n4638, n_4065);
  not g8477 (n_4066, n4650);
  and g8478 (n4651, n4638, n_4066);
  and g8479 (n4652, n_4065, n_4066);
  not g8480 (n_4067, n4651);
  not g8481 (n_4068, n4652);
  and g8482 (n4653, n_4067, n_4068);
  and g8483 (n4654, \a[1] , \a[43] );
  not g8484 (n_4069, n1367);
  not g8485 (n_4070, n4654);
  and g8486 (n4655, n_4069, n_4070);
  and g8487 (n4656, n1367, n4654);
  not g8488 (n_4071, n4655);
  not g8489 (n_4072, n4656);
  and g8490 (n4657, n_4071, n_4072);
  not g8491 (n_4073, n4657);
  and g8492 (n4658, n4431, n_4073);
  not g8493 (n_4074, n4431);
  and g8494 (n4659, n_4074, n4657);
  not g8495 (n_4075, n4658);
  not g8496 (n_4076, n4659);
  and g8497 (n4660, n_4075, n_4076);
  not g8498 (n_4077, n4415);
  and g8499 (n4661, n_4077, n4660);
  not g8500 (n_4078, n4660);
  and g8501 (n4662, n4415, n_4078);
  not g8502 (n_4079, n4661);
  not g8503 (n_4080, n4662);
  and g8504 (n4663, n_4079, n_4080);
  not g8505 (n_4081, n4653);
  and g8506 (n4664, n_4081, n4663);
  not g8507 (n_4082, n4664);
  and g8508 (n4665, n_4081, n_4082);
  and g8509 (n4666, n4663, n_4082);
  not g8510 (n_4083, n4665);
  not g8511 (n_4084, n4666);
  and g8512 (n4667, n_4083, n_4084);
  and g8513 (n4668, n_3935, n_3941);
  and g8514 (n4669, n4667, n4668);
  not g8515 (n_4085, n4667);
  not g8516 (n_4086, n4668);
  and g8517 (n4670, n_4085, n_4086);
  not g8518 (n_4087, n4669);
  not g8519 (n_4088, n4670);
  and g8520 (n4671, n_4087, n_4088);
  and g8521 (n4672, n_3918, n_3921);
  and g8522 (n4673, n_3910, n_3914);
  and g8523 (n4674, n_3786, n_3790);
  and g8524 (n4675, n4673, n4674);
  not g8525 (n_4089, n4673);
  not g8526 (n_4090, n4674);
  and g8527 (n4676, n_4089, n_4090);
  not g8528 (n_4091, n4675);
  not g8529 (n_4092, n4676);
  and g8530 (n4677, n_4091, n_4092);
  and g8531 (n4678, n_3902, n_3906);
  not g8532 (n_4093, n4677);
  and g8533 (n4679, n_4093, n4678);
  not g8534 (n_4094, n4678);
  and g8535 (n4680, n4677, n_4094);
  not g8536 (n_4095, n4679);
  not g8537 (n_4096, n4680);
  and g8538 (n4681, n_4095, n_4096);
  not g8539 (n_4097, n4672);
  and g8540 (n4682, n_4097, n4681);
  not g8541 (n_4098, n4681);
  and g8542 (n4683, n4672, n_4098);
  not g8543 (n_4099, n4682);
  not g8544 (n_4100, n4683);
  and g8545 (n4684, n_4099, n_4100);
  not g8546 (n_4101, n4671);
  not g8547 (n_4102, n4684);
  and g8548 (n4685, n_4101, n_4102);
  and g8549 (n4686, n4671, n4684);
  not g8550 (n_4103, n4686);
  and g8551 (n4687, n4635, n_4103);
  not g8552 (n_4104, n4685);
  and g8553 (n4688, n_4104, n4687);
  not g8554 (n_4105, n4688);
  and g8555 (n4689, n4635, n_4105);
  and g8556 (n4690, n_4103, n_4105);
  and g8557 (n4691, n_4104, n4690);
  not g8558 (n_4106, n4689);
  not g8559 (n_4107, n4691);
  and g8560 (n4692, n_4106, n_4107);
  and g8561 (n4693, n_3897, n_3952);
  and g8562 (n4694, n_3944, n_3948);
  and g8563 (n4695, n_3887, n_3888);
  not g8564 (n_4108, n4695);
  and g8565 (n4696, n_3893, n_4108);
  and g8566 (n4697, n4370, n4447);
  not g8567 (n_4109, n4370);
  not g8568 (n_4110, n4447);
  and g8569 (n4698, n_4109, n_4110);
  not g8570 (n_4111, n4697);
  not g8571 (n_4112, n4698);
  and g8572 (n4699, n_4111, n_4112);
  not g8573 (n_4113, n4699);
  and g8574 (n4700, n4402, n_4113);
  not g8575 (n_4114, n4402);
  and g8576 (n4701, n_4114, n4699);
  not g8577 (n_4115, n4700);
  not g8578 (n_4116, n4701);
  and g8579 (n4702, n_4115, n_4116);
  and g8580 (n4703, n_3872, n_3884);
  and g8581 (n4704, n_3835, n_3850);
  and g8582 (n4705, n4703, n4704);
  not g8583 (n_4117, n4703);
  not g8584 (n_4118, n4704);
  and g8585 (n4706, n_4117, n_4118);
  not g8586 (n_4119, n4705);
  not g8587 (n_4120, n4706);
  and g8588 (n4707, n_4119, n_4120);
  and g8589 (n4708, n4702, n4707);
  not g8590 (n_4121, n4702);
  not g8591 (n_4122, n4707);
  and g8592 (n4709, n_4121, n_4122);
  not g8593 (n_4123, n4708);
  not g8594 (n_4124, n4709);
  and g8595 (n4710, n_4123, n_4124);
  not g8596 (n_4125, n4696);
  and g8597 (n4711, n_4125, n4710);
  not g8598 (n_4126, n4710);
  and g8599 (n4712, n4696, n_4126);
  not g8600 (n_4127, n4711);
  not g8601 (n_4128, n4712);
  and g8602 (n4713, n_4127, n_4128);
  not g8603 (n_4129, n4694);
  and g8604 (n4714, n_4129, n4713);
  not g8605 (n_4130, n4713);
  and g8606 (n4715, n4694, n_4130);
  not g8607 (n_4131, n4714);
  not g8608 (n_4132, n4715);
  and g8609 (n4716, n_4131, n_4132);
  not g8610 (n_4133, n4693);
  and g8611 (n4717, n_4133, n4716);
  not g8612 (n_4134, n4716);
  and g8613 (n4718, n4693, n_4134);
  not g8614 (n_4135, n4717);
  not g8615 (n_4136, n4718);
  and g8616 (n4719, n_4135, n_4136);
  not g8617 (n_4137, n4692);
  not g8618 (n_4138, n4719);
  and g8619 (n4720, n_4137, n_4138);
  and g8620 (n4721, n4692, n4719);
  not g8621 (n_4139, n4720);
  not g8622 (n_4140, n4721);
  and g8623 (n4722, n_4139, n_4140);
  not g8624 (n_4141, n4528);
  not g8625 (n_4142, n4722);
  and g8626 (n4723, n_4141, n_4142);
  and g8627 (n4724, n4528, n4722);
  not g8628 (n_4143, n4723);
  not g8629 (n_4144, n4724);
  and g8630 (n4725, n_4143, n_4144);
  and g8631 (n4726, n_3961, n_3964);
  not g8632 (n_4145, n4726);
  and g8633 (n4727, n_3960, n_4145);
  not g8634 (n_4146, n4725);
  and g8635 (n4728, n_4146, n4727);
  not g8636 (n_4147, n4727);
  and g8637 (n4729, n4725, n_4147);
  not g8638 (n_4148, n4728);
  not g8639 (n_4149, n4729);
  and g8640 (\asquared[45] , n_4148, n_4149);
  and g8641 (n4731, n_4044, n_4047);
  and g8642 (n4732, n_4099, n_4103);
  not g8643 (n_4150, n4731);
  and g8644 (n4733, n_4150, n4732);
  not g8645 (n_4151, n4732);
  and g8646 (n4734, n4731, n_4151);
  not g8647 (n_4152, n4733);
  not g8648 (n_4153, n4734);
  and g8649 (n4735, n_4152, n_4153);
  and g8650 (n4736, n4538, n4647);
  not g8651 (n_4154, n4538);
  not g8652 (n_4155, n4647);
  and g8653 (n4737, n_4154, n_4155);
  not g8654 (n_4156, n4736);
  not g8655 (n_4157, n4737);
  and g8656 (n4738, n_4156, n_4157);
  not g8657 (n_4158, n4738);
  and g8658 (n4739, n4553, n_4158);
  not g8659 (n_4159, n4553);
  and g8660 (n4740, n_4159, n4738);
  not g8661 (n_4160, n4739);
  not g8662 (n_4161, n4740);
  and g8663 (n4741, n_4160, n_4161);
  and g8664 (n4742, n_4092, n_4096);
  not g8665 (n_4162, n4741);
  and g8666 (n4743, n_4162, n4742);
  not g8667 (n_4163, n4742);
  and g8668 (n4744, n4741, n_4163);
  not g8669 (n_4164, n4743);
  not g8670 (n_4165, n4744);
  and g8671 (n4745, n_4164, n_4165);
  and g8672 (n4746, \a[6] , \a[39] );
  not g8673 (n_4166, n3886);
  not g8674 (n_4167, n4746);
  and g8675 (n4747, n_4166, n_4167);
  and g8676 (n4748, \a[34] , \a[39] );
  and g8677 (n4749, n815, n4748);
  and g8678 (n4750, \a[12] , \a[39] );
  and g8679 (n4751, n3719, n4750);
  and g8680 (n4752, n602, n4150);
  not g8681 (n_4168, n4751);
  not g8682 (n_4169, n4752);
  and g8683 (n4753, n_4168, n_4169);
  not g8684 (n_4170, n4749);
  not g8685 (n_4171, n4753);
  and g8686 (n4754, n_4170, n_4171);
  not g8687 (n_4172, n4754);
  and g8688 (n4755, n_4170, n_4172);
  not g8689 (n_4173, n4747);
  and g8690 (n4756, n_4173, n4755);
  and g8691 (n4757, \a[33] , n_4172);
  and g8692 (n4758, \a[12] , n4757);
  not g8693 (n_4174, n4756);
  not g8694 (n_4175, n4758);
  and g8695 (n4759, n_4174, n_4175);
  and g8696 (n4760, n1048, n2334);
  and g8697 (n4761, n993, n3110);
  and g8698 (n4762, n891, n2617);
  not g8699 (n_4176, n4761);
  not g8700 (n_4177, n4762);
  and g8701 (n4763, n_4176, n_4177);
  not g8702 (n_4178, n4760);
  not g8703 (n_4179, n4763);
  and g8704 (n4764, n_4178, n_4179);
  not g8705 (n_4180, n4764);
  and g8706 (n4765, \a[30] , n_4180);
  and g8707 (n4766, \a[15] , n4765);
  and g8708 (n4767, n_4178, n_4180);
  and g8709 (n4768, \a[16] , \a[29] );
  and g8710 (n4769, \a[17] , \a[28] );
  not g8711 (n_4181, n4768);
  not g8712 (n_4182, n4769);
  and g8713 (n4770, n_4181, n_4182);
  not g8714 (n_4183, n4770);
  and g8715 (n4771, n4767, n_4183);
  not g8716 (n_4184, n4766);
  not g8717 (n_4185, n4771);
  and g8718 (n4772, n_4184, n_4185);
  not g8719 (n_4186, n4759);
  not g8720 (n_4187, n4772);
  and g8721 (n4773, n_4186, n_4187);
  not g8722 (n_4188, n4773);
  and g8723 (n4774, n_4186, n_4188);
  and g8724 (n4775, n_4187, n_4188);
  not g8725 (n_4189, n4774);
  not g8726 (n_4190, n4775);
  and g8727 (n4776, n_4189, n_4190);
  and g8728 (n4777, \a[44] , n1459);
  not g8729 (n_4191, n4777);
  and g8730 (n4778, \a[1] , n_4191);
  and g8731 (n4779, \a[44] , n4778);
  and g8732 (n4780, \a[23] , n_4191);
  not g8733 (n_4192, n4779);
  not g8734 (n_4193, n4780);
  and g8735 (n4781, n_4192, n_4193);
  and g8736 (n4782, \a[3] , \a[42] );
  not g8737 (n_4194, n4782);
  and g8738 (n4783, n_4072, n_4194);
  and g8739 (n4784, n4656, n4782);
  not g8740 (n_4195, n4781);
  not g8741 (n_4196, n4784);
  and g8742 (n4785, n_4195, n_4196);
  not g8743 (n_4197, n4783);
  and g8744 (n4786, n_4197, n4785);
  not g8745 (n_4198, n4786);
  and g8746 (n4787, n_4195, n_4198);
  and g8747 (n4788, n_4196, n_4198);
  and g8748 (n4789, n_4197, n4788);
  not g8749 (n_4199, n4787);
  not g8750 (n_4200, n4789);
  and g8751 (n4790, n_4199, n_4200);
  not g8752 (n_4201, n4776);
  not g8753 (n_4202, n4790);
  and g8754 (n4791, n_4201, n_4202);
  not g8755 (n_4203, n4791);
  and g8756 (n4792, n_4201, n_4203);
  and g8757 (n4793, n_4202, n_4203);
  not g8758 (n_4204, n4792);
  not g8759 (n_4205, n4793);
  and g8760 (n4794, n_4204, n_4205);
  not g8761 (n_4206, n4794);
  and g8762 (n4795, n4745, n_4206);
  not g8763 (n_4207, n4745);
  and g8764 (n4796, n_4207, n4794);
  not g8765 (n_4208, n4735);
  not g8766 (n_4209, n4796);
  and g8767 (n4797, n_4208, n_4209);
  not g8768 (n_4210, n4795);
  and g8769 (n4798, n_4210, n4797);
  not g8770 (n_4211, n4798);
  and g8771 (n4799, n_4208, n_4211);
  and g8772 (n4800, n_4209, n_4211);
  and g8773 (n4801, n_4210, n4800);
  not g8774 (n_4212, n4799);
  not g8775 (n_4213, n4801);
  and g8776 (n4802, n_4212, n_4213);
  and g8777 (n4803, n_4052, n_4105);
  and g8778 (n4804, n4802, n4803);
  not g8779 (n_4214, n4802);
  not g8780 (n_4215, n4803);
  and g8781 (n4805, n_4214, n_4215);
  not g8782 (n_4216, n4804);
  not g8783 (n_4217, n4805);
  and g8784 (n4806, n_4216, n_4217);
  and g8785 (n4807, \a[41] , \a[43] );
  and g8786 (n4808, n252, n4807);
  and g8787 (n4809, \a[41] , \a[45] );
  and g8788 (n4810, n212, n4809);
  and g8789 (n4811, \a[43] , \a[45] );
  and g8790 (n4812, n196, n4811);
  not g8791 (n_4219, n4810);
  not g8792 (n_4220, n4812);
  and g8793 (n4813, n_4219, n_4220);
  not g8794 (n_4221, n4808);
  not g8795 (n_4222, n4813);
  and g8796 (n4814, n_4221, n_4222);
  not g8797 (n_4223, n4814);
  and g8798 (n4815, n_4221, n_4223);
  and g8799 (n4816, \a[2] , \a[43] );
  and g8800 (n4817, \a[4] , \a[41] );
  not g8801 (n_4224, n4816);
  not g8802 (n_4225, n4817);
  and g8803 (n4818, n_4224, n_4225);
  not g8804 (n_4226, n4818);
  and g8805 (n4819, n4815, n_4226);
  and g8806 (n4820, \a[45] , n_4223);
  and g8807 (n4821, \a[0] , n4820);
  not g8808 (n_4227, n4819);
  not g8809 (n_4228, n4821);
  and g8810 (n4822, n_4227, n_4228);
  and g8811 (n4823, \a[7] , \a[38] );
  and g8812 (n4824, n432, n3687);
  and g8813 (n4825, n763, n3530);
  and g8814 (n4826, n380, n4565);
  not g8815 (n_4229, n4825);
  not g8816 (n_4230, n4826);
  and g8817 (n4827, n_4229, n_4230);
  not g8818 (n_4231, n4824);
  not g8819 (n_4232, n4827);
  and g8820 (n4828, n_4231, n_4232);
  not g8821 (n_4233, n4828);
  and g8822 (n4829, n4823, n_4233);
  and g8823 (n4830, \a[8] , \a[37] );
  and g8824 (n4831, \a[9] , \a[36] );
  not g8825 (n_4234, n4830);
  not g8826 (n_4235, n4831);
  and g8827 (n4832, n_4234, n_4235);
  and g8828 (n4833, n_4231, n_4233);
  not g8829 (n_4236, n4832);
  and g8830 (n4834, n_4236, n4833);
  not g8831 (n_4237, n4829);
  not g8832 (n_4238, n4834);
  and g8833 (n4835, n_4237, n_4238);
  not g8834 (n_4239, n4822);
  not g8835 (n_4240, n4835);
  and g8836 (n4836, n_4239, n_4240);
  not g8837 (n_4241, n4836);
  and g8838 (n4837, n_4239, n_4241);
  and g8839 (n4838, n_4240, n_4241);
  not g8840 (n_4242, n4837);
  not g8841 (n_4243, n4838);
  and g8842 (n4839, n_4242, n_4243);
  not g8843 (n_4244, n1783);
  not g8844 (n_4245, n1919);
  and g8845 (n4840, n_4244, n_4245);
  and g8846 (n4841, n1574, n1666);
  not g8847 (n_4246, n4841);
  not g8850 (n_4247, n4840);
  not g8852 (n_4248, n4844);
  and g8853 (n4845, \a[35] , n_4248);
  and g8854 (n4846, \a[10] , n4845);
  and g8855 (n4847, n_4246, n_4248);
  and g8856 (n4848, n_4247, n4847);
  not g8857 (n_4249, n4846);
  not g8858 (n_4250, n4848);
  and g8859 (n4849, n_4249, n_4250);
  not g8860 (n_4251, n4839);
  not g8861 (n_4252, n4849);
  and g8862 (n4850, n_4251, n_4252);
  not g8863 (n_4253, n4850);
  and g8864 (n4851, n_4251, n_4253);
  and g8865 (n4852, n_4252, n_4253);
  not g8866 (n_4254, n4851);
  not g8867 (n_4255, n4852);
  and g8868 (n4853, n_4254, n_4255);
  and g8869 (n4854, n745, n3812);
  and g8870 (n4855, \a[14] , \a[40] );
  and g8871 (n4856, n3100, n4855);
  not g8872 (n_4256, n4854);
  not g8873 (n_4257, n4856);
  and g8874 (n4857, n_4256, n_4257);
  and g8875 (n4858, \a[5] , \a[40] );
  and g8876 (n4859, \a[13] , \a[32] );
  and g8877 (n4860, n4858, n4859);
  not g8878 (n_4258, n4857);
  not g8879 (n_4259, n4860);
  and g8880 (n4861, n_4258, n_4259);
  not g8881 (n_4260, n4861);
  and g8882 (n4862, n_4259, n_4260);
  not g8883 (n_4261, n4858);
  not g8884 (n_4262, n4859);
  and g8885 (n4863, n_4261, n_4262);
  not g8886 (n_4263, n4863);
  and g8887 (n4864, n4862, n_4263);
  and g8888 (n4865, \a[31] , n_4260);
  and g8889 (n4866, \a[14] , n4865);
  not g8890 (n_4264, n4864);
  not g8891 (n_4265, n4866);
  and g8892 (n4867, n_4264, n_4265);
  and g8893 (n4868, n1490, n2463);
  and g8894 (n4869, n1331, n2633);
  and g8895 (n4870, n1149, n2227);
  not g8896 (n_4266, n4869);
  not g8897 (n_4267, n4870);
  and g8898 (n4871, n_4266, n_4267);
  not g8899 (n_4268, n4868);
  not g8900 (n_4269, n4871);
  and g8901 (n4872, n_4268, n_4269);
  not g8902 (n_4270, n4872);
  and g8903 (n4873, \a[27] , n_4270);
  and g8904 (n4874, \a[18] , n4873);
  and g8905 (n4875, n_4268, n_4270);
  and g8906 (n4876, \a[19] , \a[26] );
  not g8907 (n_4271, n1844);
  not g8908 (n_4272, n4876);
  and g8909 (n4877, n_4271, n_4272);
  not g8910 (n_4273, n4877);
  and g8911 (n4878, n4875, n_4273);
  not g8912 (n_4274, n4874);
  not g8913 (n_4275, n4878);
  and g8914 (n4879, n_4274, n_4275);
  not g8915 (n_4276, n4601);
  not g8916 (n_4277, n4879);
  and g8917 (n4880, n_4276, n_4277);
  not g8918 (n_4278, n4880);
  and g8919 (n4881, n_4276, n_4278);
  and g8920 (n4882, n_4277, n_4278);
  not g8921 (n_4279, n4881);
  not g8922 (n_4280, n4882);
  and g8923 (n4883, n_4279, n_4280);
  not g8924 (n_4281, n4867);
  not g8925 (n_4282, n4883);
  and g8926 (n4884, n_4281, n_4282);
  not g8927 (n_4283, n4884);
  and g8928 (n4885, n_4281, n_4283);
  and g8929 (n4886, n_4282, n_4283);
  not g8930 (n_4284, n4885);
  not g8931 (n_4285, n4886);
  and g8932 (n4887, n_4284, n_4285);
  not g8933 (n_4286, n4853);
  not g8934 (n_4287, n4887);
  and g8935 (n4888, n_4286, n_4287);
  not g8936 (n_4288, n4888);
  and g8937 (n4889, n_4286, n_4288);
  and g8938 (n4890, n_4287, n_4288);
  not g8939 (n_4289, n4889);
  not g8940 (n_4290, n4890);
  and g8941 (n4891, n_4289, n_4290);
  and g8942 (n4892, n_4120, n_4123);
  not g8943 (n_4291, n4891);
  not g8944 (n_4292, n4892);
  and g8945 (n4893, n_4291, n_4292);
  not g8946 (n_4293, n4893);
  and g8947 (n4894, n_4291, n_4293);
  and g8948 (n4895, n_4292, n_4293);
  not g8949 (n_4294, n4894);
  not g8950 (n_4295, n4895);
  and g8951 (n4896, n_4294, n_4295);
  and g8952 (n4897, n_4127, n_4131);
  and g8953 (n4898, n4896, n4897);
  not g8954 (n_4296, n4896);
  not g8955 (n_4297, n4897);
  and g8956 (n4899, n_4296, n_4297);
  not g8957 (n_4298, n4898);
  not g8958 (n_4299, n4899);
  and g8959 (n4900, n_4298, n_4299);
  and g8960 (n4901, n_4056, n_4066);
  and g8961 (n4902, n_4112, n_4116);
  and g8962 (n4903, n4901, n4902);
  not g8963 (n_4300, n4901);
  not g8964 (n_4301, n4902);
  and g8965 (n4904, n_4300, n_4301);
  not g8966 (n_4302, n4903);
  not g8967 (n_4303, n4904);
  and g8968 (n4905, n_4302, n_4303);
  and g8969 (n4906, n_4076, n_4079);
  not g8970 (n_4304, n4905);
  and g8971 (n4907, n_4304, n4906);
  not g8972 (n_4305, n4906);
  and g8973 (n4908, n4905, n_4305);
  not g8974 (n_4306, n4907);
  not g8975 (n_4307, n4908);
  and g8976 (n4909, n_4306, n_4307);
  and g8977 (n4910, n_4082, n_4088);
  not g8978 (n_4308, n4909);
  and g8979 (n4911, n_4308, n4910);
  not g8980 (n_4309, n4910);
  and g8981 (n4912, n4909, n_4309);
  not g8982 (n_4310, n4911);
  not g8983 (n_4311, n4912);
  and g8984 (n4913, n_4310, n_4311);
  and g8985 (n4914, n4570, n4587);
  not g8986 (n_4312, n4570);
  not g8987 (n_4313, n4587);
  and g8988 (n4915, n_4312, n_4313);
  not g8989 (n_4314, n4914);
  not g8990 (n_4315, n4915);
  and g8991 (n4916, n_4314, n_4315);
  not g8992 (n_4316, n4916);
  and g8993 (n4917, n4620, n_4316);
  not g8994 (n_4317, n4620);
  and g8995 (n4918, n_4317, n4916);
  not g8996 (n_4318, n4917);
  not g8997 (n_4319, n4918);
  and g8998 (n4919, n_4318, n_4319);
  and g8999 (n4920, n_4026, n_4038);
  and g9000 (n4921, n_3986, n_4001);
  and g9001 (n4922, n4920, n4921);
  not g9002 (n_4320, n4920);
  not g9003 (n_4321, n4921);
  and g9004 (n4923, n_4320, n_4321);
  not g9005 (n_4322, n4922);
  not g9006 (n_4323, n4923);
  and g9007 (n4924, n_4322, n_4323);
  and g9008 (n4925, n4919, n4924);
  not g9009 (n_4324, n4919);
  not g9010 (n_4325, n4924);
  and g9011 (n4926, n_4324, n_4325);
  not g9012 (n_4326, n4925);
  not g9013 (n_4327, n4926);
  and g9014 (n4927, n_4326, n_4327);
  and g9015 (n4928, n4913, n4927);
  not g9016 (n_4328, n4913);
  not g9017 (n_4329, n4927);
  and g9018 (n4929, n_4328, n_4329);
  not g9019 (n_4330, n4928);
  not g9020 (n_4331, n4929);
  and g9021 (n4930, n_4330, n_4331);
  and g9022 (n4931, n4900, n4930);
  not g9023 (n_4332, n4900);
  not g9024 (n_4333, n4930);
  and g9025 (n4932, n_4332, n_4333);
  not g9026 (n_4334, n4932);
  and g9027 (n4933, n4806, n_4334);
  not g9028 (n_4335, n4931);
  and g9029 (n4934, n_4335, n4933);
  not g9030 (n_4336, n4934);
  and g9031 (n4935, n4806, n_4336);
  and g9032 (n4936, n_4334, n_4336);
  and g9033 (n4937, n_4335, n4936);
  not g9034 (n_4337, n4935);
  not g9035 (n_4338, n4937);
  and g9036 (n4938, n_4337, n_4338);
  and g9037 (n4939, n_4137, n4719);
  not g9038 (n_4339, n4939);
  and g9039 (n4940, n_4135, n_4339);
  not g9040 (n_4340, n4938);
  not g9041 (n_4341, n4940);
  and g9042 (n4941, n_4340, n_4341);
  and g9043 (n4942, n4938, n4940);
  not g9044 (n_4342, n4941);
  not g9045 (n_4343, n4942);
  and g9046 (n4943, n_4342, n_4343);
  and g9047 (n4944, n_4144, n_4147);
  not g9048 (n_4344, n4944);
  and g9049 (n4945, n_4143, n_4344);
  not g9050 (n_4345, n4943);
  and g9051 (n4946, n_4345, n4945);
  not g9052 (n_4346, n4945);
  and g9053 (n4947, n4943, n_4346);
  not g9054 (n_4347, n4946);
  not g9055 (n_4348, n4947);
  and g9056 (\asquared[46] , n_4347, n_4348);
  and g9057 (n4949, n_4217, n_4336);
  and g9058 (n4950, n_4299, n_4335);
  and g9059 (n4951, n_4311, n_4330);
  and g9060 (n4952, n_4288, n_4293);
  and g9061 (n4953, n4951, n4952);
  not g9062 (n_4349, n4951);
  not g9063 (n_4350, n4952);
  and g9064 (n4954, n_4349, n_4350);
  not g9065 (n_4351, n4953);
  not g9066 (n_4352, n4954);
  and g9067 (n4955, n_4351, n_4352);
  and g9068 (n4956, \a[5] , \a[41] );
  and g9069 (n4957, \a[15] , \a[31] );
  not g9070 (n_4353, n4956);
  not g9071 (n_4354, n4957);
  and g9072 (n4958, n_4353, n_4354);
  and g9073 (n4959, \a[31] , \a[41] );
  and g9074 (n4960, n1114, n4959);
  not g9075 (n_4355, n4960);
  not g9078 (n_4356, n4958);
  not g9080 (n_4357, n4963);
  and g9081 (n4964, n_4355, n_4357);
  and g9082 (n4965, n_4356, n4964);
  and g9083 (n4966, \a[44] , n_4357);
  and g9084 (n4967, \a[2] , n4966);
  not g9085 (n_4358, n4965);
  not g9086 (n_4359, n4967);
  and g9087 (n4968, n_4358, n_4359);
  and g9088 (n4969, n745, n3143);
  and g9089 (n4970, n3419, n4855);
  not g9090 (n_4360, n4969);
  not g9091 (n_4361, n4970);
  and g9092 (n4971, n_4360, n_4361);
  and g9093 (n4972, \a[6] , \a[40] );
  and g9094 (n4973, \a[13] , \a[33] );
  and g9095 (n4974, n4972, n4973);
  not g9096 (n_4362, n4971);
  not g9097 (n_4363, n4974);
  and g9098 (n4975, n_4362, n_4363);
  not g9099 (n_4364, n4975);
  and g9100 (n4976, \a[32] , n_4364);
  and g9101 (n4977, \a[14] , n4976);
  and g9102 (n4978, n_4363, n_4364);
  not g9103 (n_4365, n4972);
  not g9104 (n_4366, n4973);
  and g9105 (n4979, n_4365, n_4366);
  not g9106 (n_4367, n4979);
  and g9107 (n4980, n4978, n_4367);
  not g9108 (n_4368, n4977);
  not g9109 (n_4369, n4980);
  and g9110 (n4981, n_4368, n_4369);
  not g9111 (n_4370, n4968);
  not g9112 (n_4371, n4981);
  and g9113 (n4982, n_4370, n_4371);
  not g9114 (n_4372, n4982);
  and g9115 (n4983, n_4370, n_4372);
  and g9116 (n4984, n_4371, n_4372);
  not g9117 (n_4373, n4983);
  not g9118 (n_4374, n4984);
  and g9119 (n4985, n_4373, n_4374);
  and g9120 (n4986, n_4315, n_4319);
  and g9121 (n4987, n4985, n4986);
  not g9122 (n_4375, n4985);
  not g9123 (n_4376, n4986);
  and g9124 (n4988, n_4375, n_4376);
  not g9125 (n_4377, n4987);
  not g9126 (n_4378, n4988);
  and g9127 (n4989, n_4377, n_4378);
  and g9128 (n4990, n4767, n4875);
  not g9129 (n_4379, n4767);
  not g9130 (n_4380, n4875);
  and g9131 (n4991, n_4379, n_4380);
  not g9132 (n_4381, n4990);
  not g9133 (n_4382, n4991);
  and g9134 (n4992, n_4381, n_4382);
  not g9135 (n_4383, n4992);
  and g9136 (n4993, n4755, n_4383);
  not g9137 (n_4384, n4755);
  and g9138 (n4994, n_4384, n4992);
  not g9139 (n_4385, n4993);
  not g9140 (n_4386, n4994);
  and g9141 (n4995, n_4385, n_4386);
  and g9142 (n4996, n_4303, n_4307);
  not g9143 (n_4387, n4995);
  and g9144 (n4997, n_4387, n4996);
  not g9145 (n_4388, n4996);
  and g9146 (n4998, n4995, n_4388);
  not g9147 (n_4389, n4997);
  not g9148 (n_4390, n4998);
  and g9149 (n4999, n_4389, n_4390);
  and g9150 (n5000, n4989, n4999);
  not g9151 (n_4391, n4989);
  not g9152 (n_4392, n4999);
  and g9153 (n5001, n_4391, n_4392);
  not g9154 (n_4393, n5000);
  not g9155 (n_4394, n5001);
  and g9156 (n5002, n_4393, n_4394);
  and g9157 (n5003, n4955, n5002);
  not g9158 (n_4395, n4955);
  not g9159 (n_4396, n5002);
  and g9160 (n5004, n_4395, n_4396);
  not g9161 (n_4397, n5003);
  not g9162 (n_4398, n5004);
  and g9163 (n5005, n_4397, n_4398);
  not g9164 (n_4399, n4950);
  and g9165 (n5006, n_4399, n5005);
  not g9166 (n_4400, n5005);
  and g9167 (n5007, n4950, n_4400);
  not g9168 (n_4401, n5006);
  not g9169 (n_4402, n5007);
  and g9170 (n5008, n_4401, n_4402);
  not g9171 (n_4403, n5008);
  and g9172 (n5009, n4949, n_4403);
  not g9173 (n_4404, n4949);
  and g9174 (n5010, n_4404, n5008);
  not g9175 (n_4405, n5009);
  not g9176 (n_4406, n5010);
  and g9177 (n5011, n_4405, n_4406);
  and g9178 (n5012, n_4150, n_4151);
  not g9179 (n_4407, n5012);
  and g9180 (n5013, n_4211, n_4407);
  and g9181 (n5014, n_4323, n_4326);
  and g9182 (n5015, \a[0] , \a[46] );
  and g9183 (n5016, \a[4] , \a[42] );
  not g9184 (n_4409, n5015);
  not g9185 (n_4410, n5016);
  and g9186 (n5017, n_4409, n_4410);
  and g9187 (n5018, \a[42] , \a[43] );
  and g9188 (n5019, n209, n5018);
  and g9189 (n5020, \a[3] , \a[46] );
  and g9190 (n5021, n4366, n5020);
  not g9191 (n_4411, n5019);
  not g9192 (n_4412, n5021);
  and g9193 (n5022, n_4411, n_4412);
  and g9194 (n5023, n5015, n5016);
  not g9195 (n_4413, n5022);
  not g9196 (n_4414, n5023);
  and g9197 (n5024, n_4413, n_4414);
  not g9198 (n_4415, n5024);
  and g9199 (n5025, n_4414, n_4415);
  not g9200 (n_4416, n5017);
  and g9201 (n5026, n_4416, n5025);
  and g9202 (n5027, \a[43] , n_4415);
  and g9203 (n5028, \a[3] , n5027);
  not g9204 (n_4417, n5026);
  not g9205 (n_4418, n5028);
  and g9206 (n5029, n_4417, n_4418);
  and g9207 (n5030, n723, n3828);
  and g9208 (n5031, \a[35] , \a[37] );
  and g9209 (n5032, n1076, n5031);
  and g9210 (n5033, n484, n3687);
  not g9211 (n_4419, n5032);
  not g9212 (n_4420, n5033);
  and g9213 (n5034, n_4419, n_4420);
  not g9214 (n_4421, n5030);
  not g9215 (n_4422, n5034);
  and g9216 (n5035, n_4421, n_4422);
  not g9217 (n_4423, n5035);
  and g9218 (n5036, \a[37] , n_4423);
  and g9219 (n5037, \a[9] , n5036);
  and g9220 (n5038, n_4421, n_4423);
  and g9221 (n5039, \a[11] , \a[35] );
  not g9222 (n_4424, n4411);
  not g9223 (n_4425, n5039);
  and g9224 (n5040, n_4424, n_4425);
  not g9225 (n_4426, n5040);
  and g9226 (n5041, n5038, n_4426);
  not g9227 (n_4427, n5037);
  not g9228 (n_4428, n5041);
  and g9229 (n5042, n_4427, n_4428);
  not g9230 (n_4429, n5029);
  not g9231 (n_4430, n5042);
  and g9232 (n5043, n_4429, n_4430);
  not g9233 (n_4431, n5043);
  and g9234 (n5044, n_4429, n_4431);
  and g9235 (n5045, n_4430, n_4431);
  not g9236 (n_4432, n5044);
  not g9237 (n_4433, n5045);
  and g9238 (n5046, n_4432, n_4433);
  and g9239 (n5047, n1494, n2463);
  and g9240 (n5048, n1492, n2633);
  and g9241 (n5049, n1490, n2227);
  not g9242 (n_4434, n5048);
  not g9243 (n_4435, n5049);
  and g9244 (n5050, n_4434, n_4435);
  not g9245 (n_4436, n5047);
  not g9246 (n_4437, n5050);
  and g9247 (n5051, n_4436, n_4437);
  not g9248 (n_4438, n5051);
  and g9249 (n5052, \a[27] , n_4438);
  and g9250 (n5053, \a[19] , n5052);
  and g9251 (n5054, n_4436, n_4438);
  and g9252 (n5055, \a[20] , \a[26] );
  and g9253 (n5056, \a[21] , \a[25] );
  not g9254 (n_4439, n5055);
  not g9255 (n_4440, n5056);
  and g9256 (n5057, n_4439, n_4440);
  not g9257 (n_4441, n5057);
  and g9258 (n5058, n5054, n_4441);
  not g9259 (n_4442, n5053);
  not g9260 (n_4443, n5058);
  and g9261 (n5059, n_4442, n_4443);
  not g9262 (n_4444, n5046);
  not g9263 (n_4445, n5059);
  and g9264 (n5060, n_4444, n_4445);
  not g9265 (n_4446, n5060);
  and g9266 (n5061, n_4444, n_4446);
  and g9267 (n5062, n_4445, n_4446);
  not g9268 (n_4447, n5061);
  not g9269 (n_4448, n5062);
  and g9270 (n5063, n_4447, n_4448);
  and g9271 (n5064, n1052, n2334);
  and g9272 (n5065, n1050, n3110);
  and g9273 (n5066, n1048, n2617);
  not g9274 (n_4449, n5065);
  not g9275 (n_4450, n5066);
  and g9276 (n5067, n_4449, n_4450);
  not g9277 (n_4451, n5064);
  not g9278 (n_4452, n5067);
  and g9279 (n5068, n_4451, n_4452);
  not g9280 (n_4453, n5068);
  and g9281 (n5069, \a[30] , n_4453);
  and g9282 (n5070, \a[16] , n5069);
  and g9283 (n5071, n_4451, n_4453);
  and g9284 (n5072, \a[17] , \a[29] );
  and g9285 (n5073, \a[18] , \a[28] );
  not g9286 (n_4454, n5072);
  not g9287 (n_4455, n5073);
  and g9288 (n5074, n_4454, n_4455);
  not g9289 (n_4456, n5074);
  and g9290 (n5075, n5071, n_4456);
  not g9291 (n_4457, n5070);
  not g9292 (n_4458, n5075);
  and g9293 (n5076, n_4457, n_4458);
  not g9294 (n_4459, n5076);
  and g9295 (n5077, n4788, n_4459);
  not g9296 (n_4460, n4788);
  and g9297 (n5078, n_4460, n5076);
  not g9298 (n_4461, n5077);
  not g9299 (n_4462, n5078);
  and g9300 (n5079, n_4461, n_4462);
  and g9301 (n5080, \a[7] , \a[39] );
  and g9302 (n5081, \a[8] , \a[38] );
  not g9303 (n_4463, n5080);
  not g9304 (n_4464, n5081);
  and g9305 (n5082, n_4463, n_4464);
  and g9306 (n5083, \a[38] , \a[39] );
  and g9307 (n5084, n380, n5083);
  not g9308 (n_4465, n5084);
  and g9309 (n5085, n3506, n_4465);
  not g9310 (n_4466, n5082);
  and g9311 (n5086, n_4466, n5085);
  not g9312 (n_4467, n5086);
  and g9313 (n5087, n3506, n_4467);
  and g9314 (n5088, n_4465, n_4467);
  and g9315 (n5089, n_4466, n5088);
  not g9316 (n_4468, n5087);
  not g9317 (n_4469, n5089);
  and g9318 (n5090, n_4468, n_4469);
  not g9319 (n_4470, n5079);
  not g9320 (n_4471, n5090);
  and g9321 (n5091, n_4470, n_4471);
  and g9322 (n5092, n5079, n5090);
  not g9323 (n_4472, n5091);
  not g9324 (n_4473, n5092);
  and g9325 (n5093, n_4472, n_4473);
  not g9326 (n_4474, n5063);
  not g9327 (n_4475, n5093);
  and g9328 (n5094, n_4474, n_4475);
  and g9329 (n5095, n5063, n5093);
  not g9330 (n_4476, n5094);
  not g9331 (n_4477, n5095);
  and g9332 (n5096, n_4476, n_4477);
  not g9333 (n_4478, n5014);
  not g9334 (n_4479, n5096);
  and g9335 (n5097, n_4478, n_4479);
  and g9336 (n5098, n5014, n5096);
  not g9337 (n_4480, n5097);
  not g9338 (n_4481, n5098);
  and g9339 (n5099, n_4480, n_4481);
  not g9340 (n_4482, n5013);
  and g9341 (n5100, n_4482, n5099);
  not g9342 (n_4483, n5099);
  and g9343 (n5101, n5013, n_4483);
  not g9344 (n_4484, n5100);
  not g9345 (n_4485, n5101);
  and g9346 (n5102, n_4484, n_4485);
  and g9347 (n5103, n_4278, n_4283);
  and g9348 (n5104, n_4241, n_4253);
  and g9349 (n5105, n5103, n5104);
  not g9350 (n_4486, n5103);
  not g9351 (n_4487, n5104);
  and g9352 (n5106, n_4486, n_4487);
  not g9353 (n_4488, n5105);
  not g9354 (n_4489, n5106);
  and g9355 (n5107, n_4488, n_4489);
  and g9356 (n5108, n_4188, n_4203);
  not g9357 (n_4490, n5107);
  and g9358 (n5109, n_4490, n5108);
  not g9359 (n_4491, n5108);
  and g9360 (n5110, n5107, n_4491);
  not g9361 (n_4492, n5109);
  not g9362 (n_4493, n5110);
  and g9363 (n5111, n_4492, n_4493);
  and g9364 (n5112, n_4165, n_4210);
  and g9365 (n5113, n4815, n4862);
  not g9366 (n_4494, n4815);
  not g9367 (n_4495, n4862);
  and g9368 (n5114, n_4494, n_4495);
  not g9369 (n_4496, n5113);
  not g9370 (n_4497, n5114);
  and g9371 (n5115, n_4496, n_4497);
  not g9372 (n_4498, n5115);
  and g9373 (n5116, n4833, n_4498);
  not g9374 (n_4499, n4833);
  and g9375 (n5117, n_4499, n5115);
  not g9376 (n_4500, n5116);
  not g9377 (n_4501, n5117);
  and g9378 (n5118, n_4500, n_4501);
  and g9379 (n5119, n_4157, n_4161);
  and g9380 (n5120, \a[1] , \a[45] );
  and g9381 (n5121, n2115, n5120);
  not g9382 (n_4502, n2115);
  not g9383 (n_4503, n5120);
  and g9384 (n5122, n_4502, n_4503);
  not g9385 (n_4504, n5121);
  not g9386 (n_4505, n5122);
  and g9387 (n5123, n_4504, n_4505);
  and g9388 (n5124, n4777, n5123);
  not g9389 (n_4506, n5124);
  and g9390 (n5125, n4777, n_4506);
  and g9391 (n5126, n_4191, n5123);
  not g9392 (n_4507, n5125);
  not g9393 (n_4508, n5126);
  and g9394 (n5127, n_4507, n_4508);
  not g9395 (n_4509, n4847);
  not g9396 (n_4510, n5127);
  and g9397 (n5128, n_4509, n_4510);
  and g9398 (n5129, n4847, n_4508);
  and g9399 (n5130, n_4507, n5129);
  not g9400 (n_4511, n5128);
  not g9401 (n_4512, n5130);
  and g9402 (n5131, n_4511, n_4512);
  not g9403 (n_4513, n5119);
  and g9404 (n5132, n_4513, n5131);
  not g9405 (n_4514, n5131);
  and g9406 (n5133, n5119, n_4514);
  not g9407 (n_4515, n5132);
  not g9408 (n_4516, n5133);
  and g9409 (n5134, n_4515, n_4516);
  and g9410 (n5135, n5118, n5134);
  not g9411 (n_4517, n5118);
  not g9412 (n_4518, n5134);
  and g9413 (n5136, n_4517, n_4518);
  not g9414 (n_4519, n5135);
  not g9415 (n_4520, n5136);
  and g9416 (n5137, n_4519, n_4520);
  not g9417 (n_4521, n5112);
  and g9418 (n5138, n_4521, n5137);
  not g9419 (n_4522, n5137);
  and g9420 (n5139, n5112, n_4522);
  not g9421 (n_4523, n5138);
  not g9422 (n_4524, n5139);
  and g9423 (n5140, n_4523, n_4524);
  and g9424 (n5141, n5111, n5140);
  not g9425 (n_4525, n5111);
  not g9426 (n_4526, n5140);
  and g9427 (n5142, n_4525, n_4526);
  not g9428 (n_4527, n5141);
  not g9429 (n_4528, n5142);
  and g9430 (n5143, n_4527, n_4528);
  and g9431 (n5144, n5102, n5143);
  not g9432 (n_4529, n5102);
  not g9433 (n_4530, n5143);
  and g9434 (n5145, n_4529, n_4530);
  not g9435 (n_4531, n5144);
  not g9436 (n_4532, n5145);
  and g9437 (n5146, n_4531, n_4532);
  not g9438 (n_4533, n5011);
  not g9439 (n_4534, n5146);
  and g9440 (n5147, n_4533, n_4534);
  and g9441 (n5148, n5011, n5146);
  not g9442 (n_4535, n5147);
  not g9443 (n_4536, n5148);
  and g9444 (n5149, n_4535, n_4536);
  and g9445 (n5150, n_4343, n_4346);
  not g9446 (n_4537, n5150);
  and g9447 (n5151, n_4342, n_4537);
  not g9448 (n_4538, n5149);
  and g9449 (n5152, n_4538, n5151);
  not g9450 (n_4539, n5151);
  and g9451 (n5153, n5149, n_4539);
  not g9452 (n_4540, n5152);
  not g9453 (n_4541, n5153);
  and g9454 (\asquared[47] , n_4540, n_4541);
  and g9455 (n5155, n_4401, n_4406);
  and g9456 (n5156, n_4352, n_4397);
  and g9457 (n5157, n_4523, n_4527);
  and g9458 (n5158, n5156, n5157);
  not g9459 (n_4542, n5156);
  not g9460 (n_4543, n5157);
  and g9461 (n5159, n_4542, n_4543);
  not g9462 (n_4544, n5158);
  not g9463 (n_4545, n5159);
  and g9464 (n5160, n_4544, n_4545);
  and g9465 (n5161, n4964, n5054);
  not g9466 (n_4546, n4964);
  not g9467 (n_4547, n5054);
  and g9468 (n5162, n_4546, n_4547);
  not g9469 (n_4548, n5161);
  not g9470 (n_4549, n5162);
  and g9471 (n5163, n_4548, n_4549);
  not g9472 (n_4550, n5163);
  and g9473 (n5164, n5025, n_4550);
  not g9474 (n_4551, n5025);
  and g9475 (n5165, n_4551, n5163);
  not g9476 (n_4552, n5164);
  not g9477 (n_4553, n5165);
  and g9478 (n5166, n_4552, n_4553);
  and g9479 (n5167, n_4431, n_4446);
  not g9480 (n_4554, n5166);
  and g9481 (n5168, n_4554, n5167);
  not g9482 (n_4555, n5167);
  and g9483 (n5169, n5166, n_4555);
  not g9484 (n_4556, n5168);
  not g9485 (n_4557, n5169);
  and g9486 (n5170, n_4556, n_4557);
  and g9487 (n5171, n_4372, n_4378);
  not g9488 (n_4558, n5170);
  and g9489 (n5172, n_4558, n5171);
  not g9490 (n_4559, n5171);
  and g9491 (n5173, n5170, n_4559);
  not g9492 (n_4560, n5172);
  not g9493 (n_4561, n5173);
  and g9494 (n5174, n_4560, n_4561);
  and g9495 (n5175, n_4474, n5093);
  not g9496 (n_4562, n5175);
  and g9497 (n5176, n_4480, n_4562);
  and g9498 (n5177, n_4390, n_4393);
  not g9499 (n_4563, n5176);
  not g9500 (n_4564, n5177);
  and g9501 (n5178, n_4563, n_4564);
  not g9502 (n_4565, n5178);
  and g9503 (n5179, n_4563, n_4565);
  and g9504 (n5180, n_4564, n_4565);
  not g9505 (n_4566, n5179);
  not g9506 (n_4567, n5180);
  and g9507 (n5181, n_4566, n_4567);
  not g9508 (n_4568, n5181);
  and g9509 (n5182, n5174, n_4568);
  not g9510 (n_4569, n5174);
  and g9511 (n5183, n_4569, n5181);
  not g9512 (n_4570, n5183);
  and g9513 (n5184, n5160, n_4570);
  not g9514 (n_4571, n5182);
  and g9515 (n5185, n_4571, n5184);
  not g9516 (n_4572, n5185);
  and g9517 (n5186, n5160, n_4572);
  and g9518 (n5187, n_4570, n_4572);
  and g9519 (n5188, n_4571, n5187);
  not g9520 (n_4573, n5186);
  not g9521 (n_4574, n5188);
  and g9522 (n5189, n_4573, n_4574);
  and g9523 (n5190, n_4484, n_4531);
  and g9524 (n5191, n_4506, n_4511);
  and g9525 (n5192, \a[12] , \a[40] );
  and g9526 (n5193, n4133, n5192);
  and g9527 (n5194, n748, n3319);
  and g9528 (n5195, \a[34] , \a[40] );
  and g9529 (n5196, n1095, n5195);
  not g9530 (n_4575, n5194);
  not g9531 (n_4576, n5196);
  and g9532 (n5197, n_4575, n_4576);
  not g9533 (n_4577, n5193);
  not g9534 (n_4578, n5197);
  and g9535 (n5198, n_4577, n_4578);
  not g9536 (n_4579, n5198);
  and g9537 (n5199, \a[34] , n_4579);
  and g9538 (n5200, \a[13] , n5199);
  and g9539 (n5201, n_4577, n_4579);
  and g9540 (n5202, \a[7] , \a[40] );
  and g9541 (n5203, \a[12] , \a[35] );
  not g9542 (n_4580, n5202);
  not g9543 (n_4581, n5203);
  and g9544 (n5204, n_4580, n_4581);
  not g9545 (n_4582, n5204);
  and g9546 (n5205, n5201, n_4582);
  not g9547 (n_4583, n5200);
  not g9548 (n_4584, n5205);
  and g9549 (n5206, n_4583, n_4584);
  not g9550 (n_4585, n5191);
  not g9551 (n_4586, n5206);
  and g9552 (n5207, n_4585, n_4586);
  not g9553 (n_4587, n5207);
  and g9554 (n5208, n_4585, n_4587);
  and g9555 (n5209, n_4586, n_4587);
  not g9556 (n_4588, n5208);
  not g9557 (n_4589, n5209);
  and g9558 (n5210, n_4588, n_4589);
  and g9559 (n5211, n_4382, n_4386);
  and g9560 (n5212, n5210, n5211);
  not g9561 (n_4590, n5210);
  not g9562 (n_4591, n5211);
  and g9563 (n5213, n_4590, n_4591);
  not g9564 (n_4592, n5212);
  not g9565 (n_4593, n5213);
  and g9566 (n5214, n_4592, n_4593);
  and g9567 (n5215, n_4515, n_4519);
  not g9568 (n_4594, n5214);
  and g9569 (n5216, n_4594, n5215);
  not g9570 (n_4595, n5215);
  and g9571 (n5217, n5214, n_4595);
  not g9572 (n_4596, n5216);
  not g9573 (n_4597, n5217);
  and g9574 (n5218, n_4596, n_4597);
  and g9575 (n5219, n_4489, n_4493);
  not g9576 (n_4598, n5218);
  and g9577 (n5220, n_4598, n5219);
  not g9578 (n_4599, n5219);
  and g9579 (n5221, n5218, n_4599);
  not g9580 (n_4600, n5220);
  not g9581 (n_4601, n5221);
  and g9582 (n5222, n_4600, n_4601);
  and g9583 (n5223, n_4460, n_4459);
  not g9584 (n_4602, n5223);
  and g9585 (n5224, n_4472, n_4602);
  and g9586 (n5225, n_4497, n_4501);
  and g9587 (n5226, n5224, n5225);
  not g9588 (n_4603, n5224);
  not g9589 (n_4604, n5225);
  and g9590 (n5227, n_4603, n_4604);
  not g9591 (n_4605, n5226);
  not g9592 (n_4606, n5227);
  and g9593 (n5228, n_4605, n_4606);
  and g9594 (n5229, \a[1] , \a[46] );
  not g9595 (n_4607, \a[24] );
  not g9596 (n_4608, n5229);
  and g9597 (n5230, n_4607, n_4608);
  and g9598 (n5231, \a[24] , \a[46] );
  and g9599 (n5232, \a[1] , n5231);
  not g9600 (n_4609, n5038);
  not g9601 (n_4610, n5232);
  and g9602 (n5233, n_4609, n_4610);
  not g9603 (n_4611, n5230);
  and g9604 (n5234, n_4611, n5233);
  not g9605 (n_4612, n5234);
  and g9606 (n5235, n_4609, n_4612);
  and g9607 (n5236, n_4610, n_4612);
  and g9608 (n5237, n_4611, n5236);
  not g9609 (n_4613, n5235);
  not g9610 (n_4614, n5237);
  and g9611 (n5238, n_4613, n_4614);
  not g9612 (n_4615, n5088);
  not g9613 (n_4616, n5238);
  and g9614 (n5239, n_4615, n_4616);
  not g9615 (n_4617, n5239);
  and g9616 (n5240, n_4615, n_4617);
  and g9617 (n5241, n_4616, n_4617);
  not g9618 (n_4618, n5240);
  not g9619 (n_4619, n5241);
  and g9620 (n5242, n_4618, n_4619);
  not g9621 (n_4620, n5242);
  and g9622 (n5243, n5228, n_4620);
  not g9623 (n_4621, n5243);
  and g9624 (n5244, n5228, n_4621);
  and g9625 (n5245, n_4620, n_4621);
  not g9626 (n_4622, n5244);
  not g9627 (n_4623, n5245);
  and g9628 (n5246, n_4622, n_4623);
  and g9629 (n5247, \a[0] , \a[47] );
  and g9630 (n5248, \a[2] , \a[45] );
  not g9631 (n_4625, n5247);
  not g9632 (n_4626, n5248);
  and g9633 (n5249, n_4625, n_4626);
  and g9634 (n5250, \a[45] , \a[47] );
  and g9635 (n5251, n196, n5250);
  not g9636 (n_4627, n5249);
  not g9637 (n_4628, n5251);
  and g9638 (n5252, n_4627, n_4628);
  and g9639 (n5253, n5121, n5252);
  not g9640 (n_4629, n5253);
  and g9641 (n5254, n_4628, n_4629);
  and g9642 (n5255, n_4627, n5254);
  and g9643 (n5256, n5121, n_4629);
  not g9644 (n_4630, n5255);
  not g9645 (n_4631, n5256);
  and g9646 (n5257, n_4630, n_4631);
  and g9647 (n5258, n1052, n2617);
  and g9648 (n5259, n1050, n3452);
  and g9649 (n5260, n1048, n2865);
  not g9650 (n_4632, n5259);
  not g9651 (n_4633, n5260);
  and g9652 (n5261, n_4632, n_4633);
  not g9653 (n_4634, n5258);
  not g9654 (n_4635, n5261);
  and g9655 (n5262, n_4634, n_4635);
  not g9656 (n_4636, n5262);
  and g9657 (n5263, \a[31] , n_4636);
  and g9658 (n5264, \a[16] , n5263);
  and g9659 (n5265, n_4634, n_4636);
  and g9660 (n5266, \a[17] , \a[30] );
  and g9661 (n5267, \a[18] , \a[29] );
  not g9662 (n_4637, n5266);
  not g9663 (n_4638, n5267);
  and g9664 (n5268, n_4637, n_4638);
  not g9665 (n_4639, n5268);
  and g9666 (n5269, n5265, n_4639);
  not g9667 (n_4640, n5264);
  not g9668 (n_4641, n5269);
  and g9669 (n5270, n_4640, n_4641);
  not g9670 (n_4642, n5257);
  not g9671 (n_4643, n5270);
  and g9672 (n5271, n_4642, n_4643);
  not g9673 (n_4644, n5271);
  and g9674 (n5272, n_4642, n_4644);
  and g9675 (n5273, n_4643, n_4644);
  not g9676 (n_4645, n5272);
  not g9677 (n_4646, n5273);
  and g9678 (n5274, n_4645, n_4646);
  and g9679 (n5275, n1494, n2227);
  and g9680 (n5276, n1492, n2800);
  and g9681 (n5277, n1490, n2331);
  not g9682 (n_4647, n5276);
  not g9683 (n_4648, n5277);
  and g9684 (n5278, n_4647, n_4648);
  not g9685 (n_4649, n5275);
  not g9686 (n_4650, n5278);
  and g9687 (n5279, n_4649, n_4650);
  not g9688 (n_4651, n5279);
  and g9689 (n5280, \a[28] , n_4651);
  and g9690 (n5281, \a[19] , n5280);
  and g9691 (n5282, n_4649, n_4651);
  and g9692 (n5283, \a[20] , \a[27] );
  not g9693 (n_4652, n2087);
  not g9694 (n_4653, n5283);
  and g9695 (n5284, n_4652, n_4653);
  not g9696 (n_4654, n5284);
  and g9697 (n5285, n5282, n_4654);
  not g9698 (n_4655, n5281);
  not g9699 (n_4656, n5285);
  and g9700 (n5286, n_4655, n_4656);
  not g9701 (n_4657, n5274);
  not g9702 (n_4658, n5286);
  and g9703 (n5287, n_4657, n_4658);
  not g9704 (n_4659, n5287);
  and g9705 (n5288, n_4657, n_4659);
  and g9706 (n5289, n_4658, n_4659);
  not g9707 (n_4660, n5288);
  not g9708 (n_4661, n5289);
  and g9709 (n5290, n_4660, n_4661);
  and g9710 (n5291, n4978, n5071);
  not g9711 (n_4662, n4978);
  not g9712 (n_4663, n5071);
  and g9713 (n5292, n_4662, n_4663);
  not g9714 (n_4664, n5291);
  not g9715 (n_4665, n5292);
  and g9716 (n5293, n_4664, n_4665);
  and g9717 (n5294, \a[32] , \a[43] );
  and g9718 (n5295, n1002, n5294);
  and g9719 (n5296, \a[43] , \a[44] );
  and g9720 (n5297, n209, n5296);
  and g9721 (n5298, \a[15] , \a[44] );
  and g9722 (n5299, n2980, n5298);
  not g9723 (n_4666, n5297);
  not g9724 (n_4667, n5299);
  and g9725 (n5300, n_4666, n_4667);
  not g9726 (n_4668, n5295);
  not g9727 (n_4669, n5300);
  and g9728 (n5301, n_4668, n_4669);
  not g9729 (n_4670, n5301);
  and g9730 (n5302, \a[44] , n_4670);
  and g9731 (n5303, \a[3] , n5302);
  and g9732 (n5304, n_4668, n_4670);
  and g9733 (n5305, \a[15] , \a[32] );
  not g9734 (n_4671, n4363);
  not g9735 (n_4672, n5305);
  and g9736 (n5306, n_4671, n_4672);
  not g9737 (n_4673, n5306);
  and g9738 (n5307, n5304, n_4673);
  not g9739 (n_4674, n5303);
  not g9740 (n_4675, n5307);
  and g9741 (n5308, n_4674, n_4675);
  not g9742 (n_4676, n5308);
  and g9743 (n5309, n5293, n_4676);
  not g9744 (n_4677, n5309);
  and g9745 (n5310, n5293, n_4677);
  and g9746 (n5311, n_4676, n_4677);
  not g9747 (n_4678, n5310);
  not g9748 (n_4679, n5311);
  and g9749 (n5312, n_4678, n_4679);
  and g9750 (n5313, n1076, n3530);
  and g9751 (n5314, n432, n5083);
  and g9752 (n5315, \a[11] , \a[39] );
  and g9753 (n5316, n4593, n5315);
  not g9754 (n_4680, n5314);
  not g9755 (n_4681, n5316);
  and g9756 (n5317, n_4680, n_4681);
  not g9757 (n_4682, n5313);
  not g9758 (n_4683, n5317);
  and g9759 (n5318, n_4682, n_4683);
  not g9760 (n_4684, n5318);
  and g9761 (n5319, n_4682, n_4684);
  and g9762 (n5320, \a[9] , \a[38] );
  and g9763 (n5321, \a[11] , \a[36] );
  not g9764 (n_4685, n5320);
  not g9765 (n_4686, n5321);
  and g9766 (n5322, n_4685, n_4686);
  not g9767 (n_4687, n5322);
  and g9768 (n5323, n5319, n_4687);
  and g9769 (n5324, \a[39] , n_4684);
  and g9770 (n5325, \a[8] , n5324);
  not g9771 (n_4688, n5323);
  not g9772 (n_4689, n5325);
  and g9773 (n5326, n_4688, n_4689);
  and g9774 (n5327, \a[22] , \a[25] );
  not g9775 (n_4690, n1666);
  not g9776 (n_4691, n5327);
  and g9777 (n5328, n_4690, n_4691);
  and g9778 (n5329, n1904, n1919);
  not g9779 (n_4692, n5329);
  not g9782 (n_4693, n5328);
  not g9784 (n_4694, n5332);
  and g9785 (n5333, \a[37] , n_4694);
  and g9786 (n5334, \a[10] , n5333);
  and g9787 (n5335, n_4692, n_4694);
  and g9788 (n5336, n_4693, n5335);
  not g9789 (n_4695, n5334);
  not g9790 (n_4696, n5336);
  and g9791 (n5337, n_4695, n_4696);
  not g9792 (n_4697, n5326);
  not g9793 (n_4698, n5337);
  and g9794 (n5338, n_4697, n_4698);
  not g9795 (n_4699, n5338);
  and g9796 (n5339, n_4697, n_4699);
  and g9797 (n5340, n_4698, n_4699);
  not g9798 (n_4700, n5339);
  not g9799 (n_4701, n5340);
  and g9800 (n5341, n_4700, n_4701);
  and g9801 (n5342, \a[33] , \a[41] );
  and g9802 (n5343, n1115, n5342);
  and g9803 (n5344, \a[41] , \a[42] );
  and g9804 (n5345, n332, n5344);
  and g9805 (n5346, \a[14] , \a[42] );
  and g9806 (n5347, n3423, n5346);
  not g9807 (n_4702, n5345);
  not g9808 (n_4703, n5347);
  and g9809 (n5348, n_4702, n_4703);
  not g9810 (n_4704, n5343);
  not g9811 (n_4705, n5348);
  and g9812 (n5349, n_4704, n_4705);
  not g9813 (n_4706, n5349);
  and g9814 (n5350, \a[42] , n_4706);
  and g9815 (n5351, \a[5] , n5350);
  and g9816 (n5352, \a[6] , \a[41] );
  and g9817 (n5353, \a[14] , \a[33] );
  not g9818 (n_4707, n5352);
  not g9819 (n_4708, n5353);
  and g9820 (n5354, n_4707, n_4708);
  and g9821 (n5355, n_4704, n_4706);
  not g9822 (n_4709, n5354);
  and g9823 (n5356, n_4709, n5355);
  not g9824 (n_4710, n5351);
  not g9825 (n_4711, n5356);
  and g9826 (n5357, n_4710, n_4711);
  not g9827 (n_4712, n5341);
  not g9828 (n_4713, n5357);
  and g9829 (n5358, n_4712, n_4713);
  not g9830 (n_4714, n5358);
  and g9831 (n5359, n_4712, n_4714);
  and g9832 (n5360, n_4713, n_4714);
  not g9833 (n_4715, n5359);
  not g9834 (n_4716, n5360);
  and g9835 (n5361, n_4715, n_4716);
  not g9836 (n_4717, n5312);
  and g9837 (n5362, n_4717, n5361);
  not g9838 (n_4718, n5361);
  and g9839 (n5363, n5312, n_4718);
  not g9840 (n_4719, n5362);
  not g9841 (n_4720, n5363);
  and g9842 (n5364, n_4719, n_4720);
  not g9843 (n_4721, n5290);
  not g9844 (n_4722, n5364);
  and g9845 (n5365, n_4721, n_4722);
  and g9846 (n5366, n5290, n5364);
  not g9847 (n_4723, n5365);
  not g9848 (n_4724, n5366);
  and g9849 (n5367, n_4723, n_4724);
  not g9850 (n_4725, n5246);
  and g9851 (n5368, n_4725, n5367);
  not g9852 (n_4726, n5368);
  and g9853 (n5369, n_4725, n_4726);
  and g9854 (n5370, n5367, n_4726);
  not g9855 (n_4727, n5369);
  not g9856 (n_4728, n5370);
  and g9857 (n5371, n_4727, n_4728);
  not g9858 (n_4729, n5371);
  and g9859 (n5372, n5222, n_4729);
  not g9860 (n_4730, n5222);
  and g9861 (n5373, n_4730, n_4728);
  and g9862 (n5374, n_4727, n5373);
  not g9863 (n_4731, n5372);
  not g9864 (n_4732, n5374);
  and g9865 (n5375, n_4731, n_4732);
  not g9866 (n_4733, n5190);
  and g9867 (n5376, n_4733, n5375);
  not g9868 (n_4734, n5376);
  and g9869 (n5377, n_4733, n_4734);
  and g9870 (n5378, n5375, n_4734);
  not g9871 (n_4735, n5377);
  not g9872 (n_4736, n5378);
  and g9873 (n5379, n_4735, n_4736);
  not g9874 (n_4737, n5189);
  not g9875 (n_4738, n5379);
  and g9876 (n5380, n_4737, n_4738);
  and g9877 (n5381, n5189, n_4736);
  and g9878 (n5382, n_4735, n5381);
  not g9879 (n_4739, n5380);
  not g9880 (n_4740, n5382);
  and g9881 (n5383, n_4739, n_4740);
  not g9882 (n_4741, n5155);
  and g9883 (n5384, n_4741, n5383);
  not g9884 (n_4742, n5383);
  and g9885 (n5385, n5155, n_4742);
  not g9886 (n_4743, n5384);
  not g9887 (n_4744, n5385);
  and g9888 (n5386, n_4743, n_4744);
  and g9889 (n5387, n_4535, n_4539);
  not g9890 (n_4745, n5387);
  and g9891 (n5388, n_4536, n_4745);
  not g9892 (n_4746, n5386);
  and g9893 (n5389, n_4746, n5388);
  not g9894 (n_4747, n5388);
  and g9895 (n5390, n5386, n_4747);
  not g9896 (n_4748, n5389);
  not g9897 (n_4749, n5390);
  and g9898 (\asquared[48] , n_4748, n_4749);
  and g9899 (n5392, n_4744, n_4747);
  not g9900 (n_4750, n5392);
  and g9901 (n5393, n_4743, n_4750);
  and g9902 (n5394, n_4734, n_4739);
  and g9903 (n5395, n_4545, n_4572);
  and g9904 (n5396, n_4565, n_4571);
  and g9905 (n5397, n_4597, n_4601);
  and g9906 (n5398, n745, n3319);
  and g9907 (n5399, n3882, n5346);
  not g9908 (n_4751, n5398);
  not g9909 (n_4752, n5399);
  and g9910 (n5400, n_4751, n_4752);
  and g9911 (n5401, \a[6] , \a[42] );
  and g9912 (n5402, \a[13] , \a[35] );
  and g9913 (n5403, n5401, n5402);
  not g9914 (n_4753, n5400);
  not g9915 (n_4754, n5403);
  and g9916 (n5404, n_4753, n_4754);
  not g9917 (n_4755, n5404);
  and g9918 (n5405, n_4754, n_4755);
  not g9919 (n_4756, n5401);
  not g9920 (n_4757, n5402);
  and g9921 (n5406, n_4756, n_4757);
  not g9922 (n_4758, n5406);
  and g9923 (n5407, n5405, n_4758);
  and g9924 (n5408, \a[34] , n_4755);
  and g9925 (n5409, \a[14] , n5408);
  not g9926 (n_4759, n5407);
  not g9927 (n_4760, n5409);
  and g9928 (n5410, n_4759, n_4760);
  and g9929 (n5411, \a[7] , \a[41] );
  and g9930 (n5412, n4593, n5192);
  and g9931 (n5413, \a[40] , \a[41] );
  and g9932 (n5414, n380, n5413);
  and g9933 (n5415, n3830, n5411);
  not g9934 (n_4761, n5414);
  not g9935 (n_4762, n5415);
  and g9936 (n5416, n_4761, n_4762);
  not g9937 (n_4763, n5412);
  not g9938 (n_4764, n5416);
  and g9939 (n5417, n_4763, n_4764);
  not g9940 (n_4765, n5417);
  and g9941 (n5418, n5411, n_4765);
  and g9942 (n5419, \a[8] , \a[40] );
  not g9943 (n_4766, n3830);
  not g9944 (n_4767, n5419);
  and g9945 (n5420, n_4766, n_4767);
  and g9946 (n5421, n_4763, n_4765);
  not g9947 (n_4768, n5420);
  and g9948 (n5422, n_4768, n5421);
  not g9949 (n_4769, n5418);
  not g9950 (n_4770, n5422);
  and g9951 (n5423, n_4769, n_4770);
  not g9952 (n_4771, n5410);
  not g9953 (n_4772, n5423);
  and g9954 (n5424, n_4771, n_4772);
  not g9955 (n_4773, n5424);
  and g9956 (n5425, n_4771, n_4773);
  and g9957 (n5426, n_4772, n_4773);
  not g9958 (n_4774, n5425);
  not g9959 (n_4775, n5426);
  and g9960 (n5427, n_4774, n_4775);
  and g9961 (n5428, \a[9] , \a[39] );
  and g9962 (n5429, n723, n4565);
  and g9963 (n5430, \a[37] , \a[39] );
  and g9964 (n5431, n1076, n5430);
  and g9965 (n5432, n484, n5083);
  not g9966 (n_4776, n5431);
  not g9967 (n_4777, n5432);
  and g9968 (n5433, n_4776, n_4777);
  not g9969 (n_4778, n5429);
  not g9970 (n_4779, n5433);
  and g9971 (n5434, n_4778, n_4779);
  not g9972 (n_4780, n5434);
  and g9973 (n5435, n5428, n_4780);
  and g9974 (n5436, n_4778, n_4780);
  and g9975 (n5437, \a[10] , \a[38] );
  not g9976 (n_4781, n4561);
  not g9977 (n_4782, n5437);
  and g9978 (n5438, n_4781, n_4782);
  not g9979 (n_4783, n5438);
  and g9980 (n5439, n5436, n_4783);
  not g9981 (n_4784, n5435);
  not g9982 (n_4785, n5439);
  and g9983 (n5440, n_4784, n_4785);
  not g9984 (n_4786, n5427);
  not g9985 (n_4787, n5440);
  and g9986 (n5441, n_4786, n_4787);
  not g9987 (n_4788, n5441);
  and g9988 (n5442, n_4786, n_4788);
  and g9989 (n5443, n_4787, n_4788);
  not g9990 (n_4789, n5442);
  not g9991 (n_4790, n5443);
  and g9992 (n5444, n_4789, n_4790);
  and g9993 (n5445, n_4587, n_4593);
  and g9994 (n5446, n5444, n5445);
  not g9995 (n_4791, n5444);
  not g9996 (n_4792, n5445);
  and g9997 (n5447, n_4791, n_4792);
  not g9998 (n_4793, n5446);
  not g9999 (n_4794, n5447);
  and g10000 (n5448, n_4793, n_4794);
  and g10001 (n5449, \a[33] , \a[43] );
  and g10002 (n5450, n1114, n5449);
  and g10003 (n5451, \a[33] , \a[44] );
  and g10004 (n5452, n1002, n5451);
  and g10005 (n5453, n226, n5296);
  not g10006 (n_4795, n5452);
  not g10007 (n_4796, n5453);
  and g10008 (n5454, n_4795, n_4796);
  not g10009 (n_4797, n5450);
  not g10010 (n_4798, n5454);
  and g10011 (n5455, n_4797, n_4798);
  not g10012 (n_4799, n5455);
  and g10013 (n5456, n_4797, n_4799);
  and g10014 (n5457, \a[5] , \a[43] );
  and g10015 (n5458, \a[15] , \a[33] );
  not g10016 (n_4800, n5457);
  not g10017 (n_4801, n5458);
  and g10018 (n5459, n_4800, n_4801);
  not g10019 (n_4802, n5459);
  and g10020 (n5460, n5456, n_4802);
  and g10021 (n5461, \a[44] , n_4799);
  and g10022 (n5462, \a[4] , n5461);
  not g10023 (n_4803, n5460);
  not g10024 (n_4804, n5462);
  and g10025 (n5463, n_4803, n_4804);
  and g10026 (n5464, n1574, n2227);
  and g10027 (n5465, n1693, n2800);
  and g10028 (n5466, n1494, n2331);
  not g10029 (n_4805, n5465);
  not g10030 (n_4806, n5466);
  and g10031 (n5467, n_4805, n_4806);
  not g10032 (n_4807, n5464);
  not g10033 (n_4808, n5467);
  and g10034 (n5468, n_4807, n_4808);
  not g10035 (n_4809, n5468);
  and g10036 (n5469, \a[28] , n_4809);
  and g10037 (n5470, \a[20] , n5469);
  and g10038 (n5471, \a[21] , \a[27] );
  and g10039 (n5472, \a[22] , \a[26] );
  not g10040 (n_4810, n5471);
  not g10041 (n_4811, n5472);
  and g10042 (n5473, n_4810, n_4811);
  and g10043 (n5474, n_4807, n_4809);
  not g10044 (n_4812, n5473);
  and g10045 (n5475, n_4812, n5474);
  not g10046 (n_4813, n5470);
  not g10047 (n_4814, n5475);
  and g10048 (n5476, n_4813, n_4814);
  not g10049 (n_4815, n5463);
  not g10050 (n_4816, n5476);
  and g10051 (n5477, n_4815, n_4816);
  not g10052 (n_4817, n5477);
  and g10053 (n5478, n_4815, n_4817);
  and g10054 (n5479, n_4816, n_4817);
  not g10055 (n_4818, n5478);
  not g10056 (n_4819, n5479);
  and g10057 (n5480, n_4818, n_4819);
  and g10058 (n5481, n1149, n2617);
  and g10059 (n5482, n3134, n3452);
  and g10060 (n5483, n1052, n2865);
  not g10061 (n_4820, n5482);
  not g10062 (n_4821, n5483);
  and g10063 (n5484, n_4820, n_4821);
  not g10064 (n_4822, n5481);
  not g10065 (n_4823, n5484);
  and g10066 (n5485, n_4822, n_4823);
  not g10067 (n_4824, n5485);
  and g10068 (n5486, \a[31] , n_4824);
  and g10069 (n5487, \a[17] , n5486);
  and g10070 (n5488, n_4822, n_4824);
  and g10071 (n5489, \a[18] , \a[30] );
  and g10072 (n5490, \a[19] , \a[29] );
  not g10073 (n_4825, n5489);
  not g10074 (n_4826, n5490);
  and g10075 (n5491, n_4825, n_4826);
  not g10076 (n_4827, n5491);
  and g10077 (n5492, n5488, n_4827);
  not g10078 (n_4828, n5487);
  not g10079 (n_4829, n5492);
  and g10080 (n5493, n_4828, n_4829);
  not g10081 (n_4830, n5480);
  not g10082 (n_4831, n5493);
  and g10083 (n5494, n_4830, n_4831);
  not g10084 (n_4832, n5494);
  and g10085 (n5495, n_4830, n_4832);
  and g10086 (n5496, n_4831, n_4832);
  not g10087 (n_4833, n5495);
  not g10088 (n_4834, n5496);
  and g10089 (n5497, n_4833, n_4834);
  not g10090 (n_4835, n5448);
  and g10091 (n5498, n_4835, n5497);
  not g10092 (n_4836, n5497);
  and g10093 (n5499, n5448, n_4836);
  not g10094 (n_4837, n5498);
  not g10095 (n_4838, n5499);
  and g10096 (n5500, n_4837, n_4838);
  not g10097 (n_4839, n5397);
  and g10098 (n5501, n_4839, n5500);
  not g10099 (n_4840, n5500);
  and g10100 (n5502, n5397, n_4840);
  not g10101 (n_4841, n5501);
  not g10102 (n_4842, n5502);
  and g10103 (n5503, n_4841, n_4842);
  not g10104 (n_4843, n5396);
  and g10105 (n5504, n_4843, n5503);
  not g10106 (n_4844, n5503);
  and g10107 (n5505, n5396, n_4844);
  not g10108 (n_4845, n5504);
  not g10109 (n_4846, n5505);
  and g10110 (n5506, n_4845, n_4846);
  not g10111 (n_4847, n5506);
  and g10112 (n5507, n5395, n_4847);
  not g10113 (n_4848, n5395);
  and g10114 (n5508, n_4848, n5506);
  not g10115 (n_4849, n5507);
  not g10116 (n_4850, n5508);
  and g10117 (n5509, n_4849, n_4850);
  and g10118 (n5510, n_4726, n_4731);
  and g10119 (n5511, n_4557, n_4561);
  and g10120 (n5512, n_4606, n_4621);
  and g10121 (n5513, n5511, n5512);
  not g10122 (n_4851, n5511);
  not g10123 (n_4852, n5512);
  and g10124 (n5514, n_4851, n_4852);
  not g10125 (n_4853, n5513);
  not g10126 (n_4854, n5514);
  and g10127 (n5515, n_4853, n_4854);
  and g10128 (n5516, \a[0] , \a[48] );
  and g10129 (n5517, n5232, n5516);
  not g10130 (n_4856, n5517);
  and g10131 (n5518, n5232, n_4856);
  and g10132 (n5519, n_4610, n5516);
  not g10133 (n_4857, n5518);
  not g10134 (n_4858, n5519);
  and g10135 (n5520, n_4857, n_4858);
  and g10136 (n5521, \a[1] , \a[47] );
  and g10137 (n5522, n1547, n5521);
  not g10138 (n_4859, n5522);
  and g10139 (n5523, n5521, n_4859);
  and g10140 (n5524, n1547, n_4859);
  not g10141 (n_4860, n5523);
  not g10142 (n_4861, n5524);
  and g10143 (n5525, n_4860, n_4861);
  not g10144 (n_4862, n5520);
  not g10145 (n_4863, n5525);
  and g10146 (n5526, n_4862, n_4863);
  not g10147 (n_4864, n5526);
  and g10148 (n5527, n_4862, n_4864);
  and g10149 (n5528, n_4863, n_4864);
  not g10150 (n_4865, n5527);
  not g10151 (n_4866, n5528);
  and g10152 (n5529, n_4865, n_4866);
  and g10153 (n5530, n_4549, n_4553);
  and g10154 (n5531, n5529, n5530);
  not g10155 (n_4867, n5529);
  not g10156 (n_4868, n5530);
  and g10157 (n5532, n_4867, n_4868);
  not g10158 (n_4869, n5531);
  not g10159 (n_4870, n5532);
  and g10160 (n5533, n_4869, n_4870);
  and g10161 (n5534, n_4665, n_4677);
  not g10162 (n_4871, n5533);
  and g10163 (n5535, n_4871, n5534);
  not g10164 (n_4872, n5534);
  and g10165 (n5536, n5533, n_4872);
  not g10166 (n_4873, n5535);
  not g10167 (n_4874, n5536);
  and g10168 (n5537, n_4873, n_4874);
  and g10169 (n5538, n5515, n5537);
  not g10170 (n_4875, n5515);
  not g10171 (n_4876, n5537);
  and g10172 (n5539, n_4875, n_4876);
  not g10173 (n_4877, n5538);
  not g10174 (n_4878, n5539);
  and g10175 (n5540, n_4877, n_4878);
  not g10176 (n_4879, n5510);
  and g10177 (n5541, n_4879, n5540);
  not g10178 (n_4880, n5541);
  and g10179 (n5542, n_4879, n_4880);
  and g10180 (n5543, n5540, n_4880);
  not g10181 (n_4881, n5542);
  not g10182 (n_4882, n5543);
  and g10183 (n5544, n_4881, n_4882);
  and g10184 (n5545, n5282, n5319);
  not g10185 (n_4883, n5282);
  not g10186 (n_4884, n5319);
  and g10187 (n5546, n_4883, n_4884);
  not g10188 (n_4885, n5545);
  not g10189 (n_4886, n5546);
  and g10190 (n5547, n_4885, n_4886);
  not g10191 (n_4887, n5547);
  and g10192 (n5548, n5355, n_4887);
  not g10193 (n_4888, n5355);
  and g10194 (n5549, n_4888, n5547);
  not g10195 (n_4889, n5548);
  not g10196 (n_4890, n5549);
  and g10197 (n5550, n_4889, n_4890);
  and g10198 (n5551, n_4699, n_4714);
  not g10199 (n_4891, n5550);
  and g10200 (n5552, n_4891, n5551);
  not g10201 (n_4892, n5551);
  and g10202 (n5553, n5550, n_4892);
  not g10203 (n_4893, n5552);
  not g10204 (n_4894, n5553);
  and g10205 (n5554, n_4893, n_4894);
  and g10206 (n5555, n5201, n5335);
  not g10207 (n_4895, n5201);
  not g10208 (n_4896, n5335);
  and g10209 (n5556, n_4895, n_4896);
  not g10210 (n_4897, n5555);
  not g10211 (n_4898, n5556);
  and g10212 (n5557, n_4897, n_4898);
  and g10213 (n5558, \a[32] , \a[46] );
  and g10214 (n5559, n902, n5558);
  and g10215 (n5560, \a[45] , \a[46] );
  and g10216 (n5561, n218, n5560);
  not g10217 (n_4899, n5559);
  not g10218 (n_4900, n5561);
  and g10219 (n5562, n_4899, n_4900);
  and g10220 (n5563, \a[3] , \a[45] );
  and g10221 (n5564, \a[16] , \a[32] );
  and g10222 (n5565, n5563, n5564);
  not g10223 (n_4901, n5562);
  not g10224 (n_4902, n5565);
  and g10225 (n5566, n_4901, n_4902);
  not g10226 (n_4903, n5566);
  and g10227 (n5567, \a[46] , n_4903);
  and g10228 (n5568, \a[2] , n5567);
  and g10229 (n5569, n_4902, n_4903);
  not g10230 (n_4904, n5563);
  not g10231 (n_4905, n5564);
  and g10232 (n5570, n_4904, n_4905);
  not g10233 (n_4906, n5570);
  and g10234 (n5571, n5569, n_4906);
  not g10235 (n_4907, n5568);
  not g10236 (n_4908, n5571);
  and g10237 (n5572, n_4907, n_4908);
  not g10238 (n_4909, n5572);
  and g10239 (n5573, n5557, n_4909);
  not g10240 (n_4910, n5573);
  and g10241 (n5574, n5557, n_4910);
  and g10242 (n5575, n_4909, n_4910);
  not g10243 (n_4911, n5574);
  not g10244 (n_4912, n5575);
  and g10245 (n5576, n_4911, n_4912);
  not g10246 (n_4913, n5554);
  and g10247 (n5577, n_4913, n5576);
  not g10248 (n_4914, n5576);
  and g10249 (n5578, n5554, n_4914);
  not g10250 (n_4915, n5577);
  not g10251 (n_4916, n5578);
  and g10252 (n5579, n_4915, n_4916);
  and g10253 (n5580, n_4717, n_4718);
  not g10254 (n_4917, n5580);
  and g10255 (n5581, n_4723, n_4917);
  not g10256 (n_4918, n5581);
  and g10257 (n5582, n5579, n_4918);
  not g10258 (n_4919, n5579);
  and g10259 (n5583, n_4919, n5581);
  not g10260 (n_4920, n5582);
  not g10261 (n_4921, n5583);
  and g10262 (n5584, n_4920, n_4921);
  and g10263 (n5585, n5265, n5304);
  not g10264 (n_4922, n5265);
  not g10265 (n_4923, n5304);
  and g10266 (n5586, n_4922, n_4923);
  not g10267 (n_4924, n5585);
  not g10268 (n_4925, n5586);
  and g10269 (n5587, n_4924, n_4925);
  not g10270 (n_4926, n5587);
  and g10271 (n5588, n5254, n_4926);
  not g10272 (n_4927, n5254);
  and g10273 (n5589, n_4927, n5587);
  not g10274 (n_4928, n5588);
  not g10275 (n_4929, n5589);
  and g10276 (n5590, n_4928, n_4929);
  and g10277 (n5591, n_4612, n_4617);
  and g10278 (n5592, n_4644, n_4659);
  and g10279 (n5593, n5591, n5592);
  not g10280 (n_4930, n5591);
  not g10281 (n_4931, n5592);
  and g10282 (n5594, n_4930, n_4931);
  not g10283 (n_4932, n5593);
  not g10284 (n_4933, n5594);
  and g10285 (n5595, n_4932, n_4933);
  and g10286 (n5596, n5590, n5595);
  not g10287 (n_4934, n5590);
  not g10288 (n_4935, n5595);
  and g10289 (n5597, n_4934, n_4935);
  not g10290 (n_4936, n5596);
  not g10291 (n_4937, n5597);
  and g10292 (n5598, n_4936, n_4937);
  and g10293 (n5599, n5584, n5598);
  not g10294 (n_4938, n5584);
  not g10295 (n_4939, n5598);
  and g10296 (n5600, n_4938, n_4939);
  not g10297 (n_4940, n5599);
  not g10298 (n_4941, n5600);
  and g10299 (n5601, n_4940, n_4941);
  not g10300 (n_4942, n5544);
  and g10301 (n5602, n_4942, n5601);
  not g10302 (n_4943, n5601);
  and g10303 (n5603, n_4882, n_4943);
  and g10304 (n5604, n_4881, n5603);
  not g10305 (n_4944, n5602);
  not g10306 (n_4945, n5604);
  and g10307 (n5605, n_4944, n_4945);
  and g10308 (n5606, n5509, n5605);
  not g10309 (n_4946, n5509);
  not g10310 (n_4947, n5605);
  and g10311 (n5607, n_4946, n_4947);
  not g10312 (n_4948, n5606);
  not g10313 (n_4949, n5607);
  and g10314 (n5608, n_4948, n_4949);
  not g10315 (n_4950, n5608);
  and g10316 (n5609, n5394, n_4950);
  not g10317 (n_4951, n5394);
  and g10318 (n5610, n_4951, n5608);
  not g10319 (n_4952, n5609);
  not g10320 (n_4953, n5610);
  and g10321 (n5611, n_4952, n_4953);
  not g10322 (n_4954, n5611);
  and g10323 (n5612, n5393, n_4954);
  not g10324 (n_4955, n5393);
  and g10325 (n5613, n_4955, n_4952);
  and g10326 (n5614, n_4953, n5613);
  not g10327 (n_4956, n5612);
  not g10328 (n_4957, n5614);
  and g10329 (\asquared[49] , n_4956, n_4957);
  and g10330 (n5616, n_4880, n_4944);
  and g10331 (n5617, n_4920, n_4940);
  and g10332 (n5618, n_4854, n_4877);
  and g10333 (n5619, \a[7] , \a[42] );
  and g10334 (n5620, \a[8] , \a[41] );
  not g10335 (n_4958, n5619);
  not g10336 (n_4959, n5620);
  and g10337 (n5621, n_4958, n_4959);
  and g10338 (n5622, n380, n5344);
  not g10339 (n_4960, n5622);
  not g10342 (n_4961, n5621);
  not g10344 (n_4962, n5625);
  and g10345 (n5626, n_4960, n_4962);
  and g10346 (n5627, n_4961, n5626);
  and g10347 (n5628, \a[36] , n_4962);
  and g10348 (n5629, \a[13] , n5628);
  not g10349 (n_4963, n5627);
  not g10350 (n_4964, n5629);
  and g10351 (n5630, n_4963, n_4964);
  not g10352 (n_4965, n1904);
  not g10353 (n_4966, n2303);
  and g10354 (n5631, n_4965, n_4966);
  and g10355 (n5632, n1904, n2303);
  not g10356 (n_4967, n5632);
  not g10359 (n_4968, n5631);
  not g10361 (n_4969, n5635);
  and g10362 (n5636, \a[38] , n_4969);
  and g10363 (n5637, \a[11] , n5636);
  and g10364 (n5638, n_4967, n_4969);
  and g10365 (n5639, n_4968, n5638);
  not g10366 (n_4970, n5637);
  not g10367 (n_4971, n5639);
  and g10368 (n5640, n_4970, n_4971);
  not g10369 (n_4972, n5630);
  not g10370 (n_4973, n5640);
  and g10371 (n5641, n_4972, n_4973);
  not g10372 (n_4974, n5641);
  and g10373 (n5642, n_4972, n_4974);
  and g10374 (n5643, n_4973, n_4974);
  not g10375 (n_4975, n5642);
  not g10376 (n_4976, n5643);
  and g10377 (n5644, n_4975, n_4976);
  and g10378 (n5645, \a[35] , \a[43] );
  and g10379 (n5646, n1115, n5645);
  and g10380 (n5647, \a[15] , \a[43] );
  and g10381 (n5648, n3882, n5647);
  and g10382 (n5649, n895, n3319);
  not g10383 (n_4977, n5648);
  not g10384 (n_4978, n5649);
  and g10385 (n5650, n_4977, n_4978);
  not g10386 (n_4979, n5646);
  not g10387 (n_4980, n5650);
  and g10388 (n5651, n_4979, n_4980);
  not g10389 (n_4981, n5651);
  and g10390 (n5652, \a[34] , n_4981);
  and g10391 (n5653, \a[15] , n5652);
  and g10392 (n5654, \a[6] , \a[43] );
  and g10393 (n5655, \a[14] , \a[35] );
  not g10394 (n_4982, n5654);
  not g10395 (n_4983, n5655);
  and g10396 (n5656, n_4982, n_4983);
  and g10397 (n5657, n_4979, n_4981);
  not g10398 (n_4984, n5656);
  and g10399 (n5658, n_4984, n5657);
  not g10400 (n_4985, n5653);
  not g10401 (n_4986, n5658);
  and g10402 (n5659, n_4985, n_4986);
  not g10403 (n_4987, n5644);
  not g10404 (n_4988, n5659);
  and g10405 (n5660, n_4987, n_4988);
  not g10406 (n_4989, n5660);
  and g10407 (n5661, n_4987, n_4989);
  and g10408 (n5662, n_4988, n_4989);
  not g10409 (n_4990, n5661);
  not g10410 (n_4991, n5662);
  and g10411 (n5663, n_4990, n_4991);
  and g10412 (n5664, \a[2] , \a[47] );
  not g10413 (n_4992, n5020);
  not g10414 (n_4993, n5664);
  and g10415 (n5665, n_4992, n_4993);
  and g10416 (n5666, \a[46] , \a[47] );
  and g10417 (n5667, n218, n5666);
  not g10418 (n_4994, n5667);
  not g10421 (n_4995, n5665);
  not g10423 (n_4996, n5670);
  and g10424 (n5671, n_4994, n_4996);
  and g10425 (n5672, n_4995, n5671);
  and g10426 (n5673, \a[27] , n_4996);
  and g10427 (n5674, \a[22] , n5673);
  not g10428 (n_4997, n5672);
  not g10429 (n_4998, n5674);
  and g10430 (n5675, n_4997, n_4998);
  and g10431 (n5676, n1494, n2334);
  and g10432 (n5677, n1492, n3110);
  and g10433 (n5678, n1490, n2617);
  not g10434 (n_4999, n5677);
  not g10435 (n_5000, n5678);
  and g10436 (n5679, n_4999, n_5000);
  not g10437 (n_5001, n5676);
  not g10438 (n_5002, n5679);
  and g10439 (n5680, n_5001, n_5002);
  not g10440 (n_5003, n5680);
  and g10441 (n5681, \a[30] , n_5003);
  and g10442 (n5682, \a[19] , n5681);
  and g10443 (n5683, n_5001, n_5003);
  and g10444 (n5684, \a[20] , \a[29] );
  and g10445 (n5685, \a[21] , \a[28] );
  not g10446 (n_5004, n5684);
  not g10447 (n_5005, n5685);
  and g10448 (n5686, n_5004, n_5005);
  not g10449 (n_5006, n5686);
  and g10450 (n5687, n5683, n_5006);
  not g10451 (n_5007, n5682);
  not g10452 (n_5008, n5687);
  and g10453 (n5688, n_5007, n_5008);
  not g10454 (n_5009, n5675);
  not g10455 (n_5010, n5688);
  and g10456 (n5689, n_5009, n_5010);
  not g10457 (n_5011, n5689);
  and g10458 (n5690, n_5009, n_5011);
  and g10459 (n5691, n_5010, n_5011);
  not g10460 (n_5012, n5690);
  not g10461 (n_5013, n5691);
  and g10462 (n5692, n_5012, n_5013);
  and g10463 (n5693, n480, n5430);
  and g10464 (n5694, n484, n4171);
  and g10465 (n5695, \a[37] , \a[40] );
  and g10466 (n5696, n1182, n5695);
  not g10467 (n_5014, n5694);
  not g10468 (n_5015, n5696);
  and g10469 (n5697, n_5014, n_5015);
  not g10470 (n_5016, n5693);
  not g10471 (n_5017, n5697);
  and g10472 (n5698, n_5016, n_5017);
  not g10473 (n_5018, n5698);
  and g10474 (n5699, \a[40] , n_5018);
  and g10475 (n5700, \a[9] , n5699);
  and g10476 (n5701, n_5016, n_5018);
  and g10477 (n5702, \a[10] , \a[39] );
  not g10478 (n_5019, n4485);
  not g10479 (n_5020, n5702);
  and g10480 (n5703, n_5019, n_5020);
  not g10481 (n_5021, n5703);
  and g10482 (n5704, n5701, n_5021);
  not g10483 (n_5022, n5700);
  not g10484 (n_5023, n5704);
  and g10485 (n5705, n_5022, n_5023);
  not g10486 (n_5024, n5692);
  not g10487 (n_5025, n5705);
  and g10488 (n5706, n_5024, n_5025);
  not g10489 (n_5026, n5706);
  and g10490 (n5707, n_5024, n_5026);
  and g10491 (n5708, n_5025, n_5026);
  not g10492 (n_5027, n5707);
  not g10493 (n_5028, n5708);
  and g10494 (n5709, n_5027, n_5028);
  and g10495 (n5710, \a[44] , n224);
  and g10496 (n5711, \a[45] , n212);
  not g10497 (n_5029, n5710);
  not g10498 (n_5030, n5711);
  and g10499 (n5712, n_5029, n_5030);
  and g10500 (n5713, \a[44] , \a[45] );
  and g10501 (n5714, n226, n5713);
  not g10502 (n_5032, n5714);
  and g10503 (n5715, \a[49] , n_5032);
  not g10504 (n_5033, n5712);
  and g10505 (n5716, n_5033, n5715);
  not g10506 (n_5034, n5716);
  and g10507 (n5717, \a[0] , n_5034);
  and g10508 (n5718, \a[49] , n5717);
  and g10509 (n5719, n_5032, n_5034);
  and g10510 (n5720, \a[4] , \a[45] );
  and g10511 (n5721, \a[5] , \a[44] );
  not g10512 (n_5035, n5720);
  not g10513 (n_5036, n5721);
  and g10514 (n5722, n_5035, n_5036);
  not g10515 (n_5037, n5722);
  and g10516 (n5723, n5719, n_5037);
  not g10517 (n_5038, n5718);
  not g10518 (n_5039, n5723);
  and g10519 (n5724, n_5038, n_5039);
  and g10520 (n5725, n_4856, n_4864);
  not g10521 (n_5040, n5724);
  and g10522 (n5726, n_5040, n5725);
  not g10523 (n_5041, n5725);
  and g10524 (n5727, n5724, n_5041);
  not g10525 (n_5042, n5726);
  not g10526 (n_5043, n5727);
  and g10527 (n5728, n_5042, n_5043);
  and g10528 (n5729, n1052, n3812);
  and g10529 (n5730, n1050, n2598);
  and g10530 (n5731, n1048, n3143);
  not g10531 (n_5044, n5730);
  not g10532 (n_5045, n5731);
  and g10533 (n5732, n_5044, n_5045);
  not g10534 (n_5046, n5729);
  not g10535 (n_5047, n5732);
  and g10536 (n5733, n_5046, n_5047);
  not g10537 (n_5048, n5733);
  and g10538 (n5734, \a[33] , n_5048);
  and g10539 (n5735, \a[16] , n5734);
  and g10540 (n5736, n_5046, n_5048);
  and g10541 (n5737, \a[17] , \a[32] );
  and g10542 (n5738, \a[18] , \a[31] );
  not g10543 (n_5049, n5737);
  not g10544 (n_5050, n5738);
  and g10545 (n5739, n_5049, n_5050);
  not g10546 (n_5051, n5739);
  and g10547 (n5740, n5736, n_5051);
  not g10548 (n_5052, n5735);
  not g10549 (n_5053, n5740);
  and g10550 (n5741, n_5052, n_5053);
  not g10551 (n_5054, n5728);
  not g10552 (n_5055, n5741);
  and g10553 (n5742, n_5054, n_5055);
  and g10554 (n5743, n5728, n5741);
  not g10555 (n_5056, n5742);
  not g10556 (n_5057, n5743);
  and g10557 (n5744, n_5056, n_5057);
  and g10558 (n5745, n5709, n5744);
  not g10559 (n_5058, n5709);
  not g10560 (n_5059, n5744);
  and g10561 (n5746, n_5058, n_5059);
  not g10562 (n_5060, n5745);
  not g10563 (n_5061, n5746);
  and g10564 (n5747, n_5060, n_5061);
  not g10565 (n_5062, n5663);
  not g10566 (n_5063, n5747);
  and g10567 (n5748, n_5062, n_5063);
  and g10568 (n5749, n5663, n5747);
  not g10569 (n_5064, n5748);
  not g10570 (n_5065, n5749);
  and g10571 (n5750, n_5064, n_5065);
  not g10572 (n_5066, n5618);
  and g10573 (n5751, n_5066, n5750);
  not g10574 (n_5067, n5750);
  and g10575 (n5752, n5618, n_5067);
  not g10576 (n_5068, n5751);
  not g10577 (n_5069, n5752);
  and g10578 (n5753, n_5068, n_5069);
  not g10579 (n_5070, n5617);
  and g10580 (n5754, n_5070, n5753);
  not g10581 (n_5071, n5753);
  and g10582 (n5755, n5617, n_5071);
  not g10583 (n_5072, n5754);
  not g10584 (n_5073, n5755);
  and g10585 (n5756, n_5072, n_5073);
  not g10586 (n_5074, n5616);
  and g10587 (n5757, n_5074, n5756);
  not g10588 (n_5075, n5756);
  and g10589 (n5758, n5616, n_5075);
  not g10590 (n_5076, n5757);
  not g10591 (n_5077, n5758);
  and g10592 (n5759, n_5076, n_5077);
  and g10593 (n5760, n_4841, n_4845);
  and g10594 (n5761, n_4886, n_4890);
  and g10595 (n5762, n_4898, n_4910);
  and g10596 (n5763, n5761, n5762);
  not g10597 (n_5078, n5761);
  not g10598 (n_5079, n5762);
  and g10599 (n5764, n_5078, n_5079);
  not g10600 (n_5080, n5763);
  not g10601 (n_5081, n5764);
  and g10602 (n5765, n_5080, n_5081);
  and g10603 (n5766, n_4925, n_4929);
  not g10604 (n_5082, n5765);
  and g10605 (n5767, n_5082, n5766);
  not g10606 (n_5083, n5766);
  and g10607 (n5768, n5765, n_5083);
  not g10608 (n_5084, n5767);
  not g10609 (n_5085, n5768);
  and g10610 (n5769, n_5084, n_5085);
  and g10611 (n5770, n_4894, n_4916);
  and g10612 (n5771, n_4933, n_4936);
  not g10613 (n_5086, n5770);
  not g10614 (n_5087, n5771);
  and g10615 (n5772, n_5086, n_5087);
  not g10616 (n_5088, n5772);
  and g10617 (n5773, n_5086, n_5088);
  and g10618 (n5774, n_5087, n_5088);
  not g10619 (n_5089, n5773);
  not g10620 (n_5090, n5774);
  and g10621 (n5775, n_5089, n_5090);
  not g10622 (n_5091, n5769);
  and g10623 (n5776, n_5091, n5775);
  not g10624 (n_5092, n5775);
  and g10625 (n5777, n5769, n_5092);
  not g10626 (n_5093, n5776);
  not g10627 (n_5094, n5777);
  and g10628 (n5778, n_5093, n_5094);
  not g10629 (n_5095, n5760);
  and g10630 (n5779, n_5095, n5778);
  not g10631 (n_5096, n5779);
  and g10632 (n5780, n_5095, n_5096);
  and g10633 (n5781, n5778, n_5096);
  not g10634 (n_5097, n5780);
  not g10635 (n_5098, n5781);
  and g10636 (n5782, n_5097, n_5098);
  and g10637 (n5783, n5405, n5488);
  not g10638 (n_5099, n5405);
  not g10639 (n_5100, n5488);
  and g10640 (n5784, n_5099, n_5100);
  not g10641 (n_5101, n5783);
  not g10642 (n_5102, n5784);
  and g10643 (n5785, n_5101, n_5102);
  not g10644 (n_5103, n5785);
  and g10645 (n5786, n5421, n_5103);
  not g10646 (n_5104, n5421);
  and g10647 (n5787, n_5104, n5785);
  not g10648 (n_5105, n5786);
  not g10649 (n_5106, n5787);
  and g10650 (n5788, n_5105, n_5106);
  and g10651 (n5789, n_4817, n_4832);
  not g10652 (n_5107, n5788);
  and g10653 (n5790, n_5107, n5789);
  not g10654 (n_5108, n5789);
  and g10655 (n5791, n5788, n_5108);
  not g10656 (n_5109, n5790);
  not g10657 (n_5110, n5791);
  and g10658 (n5792, n_5109, n_5110);
  and g10659 (n5793, n_4870, n_4874);
  not g10660 (n_5111, n5792);
  and g10661 (n5794, n_5111, n5793);
  not g10662 (n_5112, n5793);
  and g10663 (n5795, n5792, n_5112);
  not g10664 (n_5113, n5794);
  not g10665 (n_5114, n5795);
  and g10666 (n5796, n_5113, n_5114);
  and g10667 (n5797, n_4794, n_4838);
  not g10668 (n_5115, n5797);
  and g10669 (n5798, n5796, n_5115);
  not g10670 (n_5116, n5796);
  and g10671 (n5799, n_5116, n5797);
  not g10672 (n_5117, n5798);
  not g10673 (n_5118, n5799);
  and g10674 (n5800, n_5117, n_5118);
  and g10675 (n5801, n5456, n5569);
  not g10676 (n_5119, n5456);
  not g10677 (n_5120, n5569);
  and g10678 (n5802, n_5119, n_5120);
  not g10679 (n_5121, n5801);
  not g10680 (n_5122, n5802);
  and g10681 (n5803, n_5121, n_5122);
  not g10682 (n_5123, n5803);
  and g10683 (n5804, n5474, n_5123);
  not g10684 (n_5124, n5474);
  and g10685 (n5805, n_5124, n5803);
  not g10686 (n_5125, n5804);
  not g10687 (n_5126, n5805);
  and g10688 (n5806, n_5125, n_5126);
  and g10689 (n5807, n_4773, n_4788);
  and g10690 (n5808, \a[48] , n1747);
  and g10691 (n5809, \a[1] , \a[48] );
  not g10692 (n_5127, \a[25] );
  not g10693 (n_5128, n5809);
  and g10694 (n5810, n_5127, n_5128);
  not g10695 (n_5129, n5808);
  not g10696 (n_5130, n5810);
  and g10697 (n5811, n_5129, n_5130);
  and g10698 (n5812, n5522, n5811);
  not g10699 (n_5131, n5811);
  and g10700 (n5813, n_4859, n_5131);
  not g10701 (n_5132, n5812);
  not g10702 (n_5133, n5813);
  and g10703 (n5814, n_5132, n_5133);
  not g10704 (n_5134, n5436);
  and g10705 (n5815, n_5134, n5814);
  not g10706 (n_5135, n5814);
  and g10707 (n5816, n5436, n_5135);
  not g10708 (n_5136, n5815);
  not g10709 (n_5137, n5816);
  and g10710 (n5817, n_5136, n_5137);
  not g10711 (n_5138, n5807);
  and g10712 (n5818, n_5138, n5817);
  not g10713 (n_5139, n5817);
  and g10714 (n5819, n5807, n_5139);
  not g10715 (n_5140, n5818);
  not g10716 (n_5141, n5819);
  and g10717 (n5820, n_5140, n_5141);
  and g10718 (n5821, n5806, n5820);
  not g10719 (n_5142, n5806);
  not g10720 (n_5143, n5820);
  and g10721 (n5822, n_5142, n_5143);
  not g10722 (n_5144, n5821);
  not g10723 (n_5145, n5822);
  and g10724 (n5823, n_5144, n_5145);
  and g10725 (n5824, n5800, n5823);
  not g10726 (n_5146, n5800);
  not g10727 (n_5147, n5823);
  and g10728 (n5825, n_5146, n_5147);
  not g10729 (n_5148, n5824);
  not g10730 (n_5149, n5825);
  and g10731 (n5826, n_5148, n_5149);
  not g10732 (n_5150, n5782);
  and g10733 (n5827, n_5150, n5826);
  not g10734 (n_5151, n5826);
  and g10735 (n5828, n_5098, n_5151);
  and g10736 (n5829, n_5097, n5828);
  not g10737 (n_5152, n5827);
  not g10738 (n_5153, n5829);
  and g10739 (n5830, n_5152, n_5153);
  and g10740 (n5831, n5759, n5830);
  not g10741 (n_5154, n5759);
  not g10742 (n_5155, n5830);
  and g10743 (n5832, n_5154, n_5155);
  not g10744 (n_5156, n5831);
  not g10745 (n_5157, n5832);
  and g10746 (n5833, n_5156, n_5157);
  and g10747 (n5834, n_4850, n_4948);
  not g10748 (n_5158, n5833);
  and g10749 (n5835, n_5158, n5834);
  not g10750 (n_5159, n5834);
  and g10751 (n5836, n5833, n_5159);
  not g10752 (n_5160, n5835);
  not g10753 (n_5161, n5836);
  and g10754 (n5837, n_5160, n_5161);
  not g10755 (n_5162, n5613);
  and g10756 (n5838, n_4953, n_5162);
  not g10757 (n_5163, n5837);
  and g10758 (n5839, n_5163, n5838);
  not g10759 (n_5164, n5838);
  and g10760 (n5840, n5837, n_5164);
  not g10761 (n_5165, n5839);
  not g10762 (n_5166, n5840);
  and g10763 (\asquared[50] , n_5165, n_5166);
  and g10764 (n5842, n_5160, n_5164);
  not g10765 (n_5167, n5842);
  and g10766 (n5843, n_5161, n_5167);
  and g10767 (n5844, n_5076, n_5156);
  and g10768 (n5845, n_5096, n_5152);
  and g10769 (n5846, n_5117, n_5148);
  and g10770 (n5847, n_5088, n_5094);
  and g10771 (n5848, \a[35] , \a[45] );
  and g10772 (n5849, n1114, n5848);
  and g10773 (n5850, \a[16] , \a[45] );
  and g10774 (n5851, n3664, n5850);
  and g10775 (n5852, n891, n3319);
  not g10776 (n_5168, n5851);
  not g10777 (n_5169, n5852);
  and g10778 (n5853, n_5168, n_5169);
  not g10779 (n_5170, n5849);
  not g10780 (n_5171, n5853);
  and g10781 (n5854, n_5170, n_5171);
  not g10782 (n_5172, n5854);
  and g10783 (n5855, n_5170, n_5172);
  and g10784 (n5856, \a[5] , \a[45] );
  and g10785 (n5857, \a[15] , \a[35] );
  not g10786 (n_5173, n5856);
  not g10787 (n_5174, n5857);
  and g10788 (n5858, n_5173, n_5174);
  not g10789 (n_5175, n5858);
  and g10790 (n5859, n5855, n_5175);
  and g10791 (n5860, \a[34] , n_5172);
  and g10792 (n5861, \a[16] , n5860);
  not g10793 (n_5176, n5859);
  not g10794 (n_5177, n5861);
  and g10795 (n5862, n_5176, n_5177);
  and g10796 (n5863, \a[28] , \a[32] );
  and g10797 (n5864, n1469, n5863);
  and g10798 (n5865, n1919, n2331);
  not g10799 (n_5178, n5864);
  not g10800 (n_5179, n5865);
  and g10801 (n5866, n_5178, n_5179);
  and g10802 (n5867, \a[18] , \a[32] );
  and g10803 (n5868, \a[23] , \a[27] );
  and g10804 (n5869, n5867, n5868);
  not g10805 (n_5180, n5866);
  not g10806 (n_5181, n5869);
  and g10807 (n5870, n_5180, n_5181);
  not g10808 (n_5182, n5870);
  and g10809 (n5871, \a[28] , n_5182);
  and g10810 (n5872, \a[22] , n5871);
  not g10811 (n_5183, n5867);
  not g10812 (n_5184, n5868);
  and g10813 (n5873, n_5183, n_5184);
  and g10814 (n5874, n_5181, n_5182);
  not g10815 (n_5185, n5873);
  and g10816 (n5875, n_5185, n5874);
  not g10817 (n_5186, n5872);
  not g10818 (n_5187, n5875);
  and g10819 (n5876, n_5186, n_5187);
  not g10820 (n_5188, n5862);
  not g10821 (n_5189, n5876);
  and g10822 (n5877, n_5188, n_5189);
  not g10823 (n_5190, n5877);
  and g10824 (n5878, n_5188, n_5190);
  and g10825 (n5879, n_5189, n_5190);
  not g10826 (n_5191, n5878);
  not g10827 (n_5192, n5879);
  and g10828 (n5880, n_5191, n_5192);
  and g10829 (n5881, n_5132, n_5136);
  and g10830 (n5882, n5880, n5881);
  not g10831 (n_5193, n5880);
  not g10832 (n_5194, n5881);
  and g10833 (n5883, n_5193, n_5194);
  not g10834 (n_5195, n5882);
  not g10835 (n_5196, n5883);
  and g10836 (n5884, n_5195, n_5196);
  and g10837 (n5885, \a[0] , \a[50] );
  and g10838 (n5886, \a[2] , \a[48] );
  not g10839 (n_5198, n5885);
  not g10840 (n_5199, n5886);
  and g10841 (n5887, n_5198, n_5199);
  and g10842 (n5888, \a[48] , \a[50] );
  and g10843 (n5889, n196, n5888);
  not g10844 (n_5200, n5887);
  not g10845 (n_5201, n5889);
  and g10846 (n5890, n_5200, n_5201);
  and g10847 (n5891, n5808, n5890);
  not g10848 (n_5202, n5891);
  and g10849 (n5892, n_5201, n_5202);
  and g10850 (n5893, n_5200, n5892);
  and g10851 (n5894, n5808, n_5202);
  not g10852 (n_5203, n5893);
  not g10853 (n_5204, n5894);
  and g10854 (n5895, n_5203, n_5204);
  and g10855 (n5896, \a[33] , \a[46] );
  and g10856 (n5897, n1181, n5896);
  and g10857 (n5898, n209, n5666);
  and g10858 (n5899, \a[17] , \a[47] );
  and g10859 (n5900, n3146, n5899);
  not g10860 (n_5205, n5898);
  not g10861 (n_5206, n5900);
  and g10862 (n5901, n_5205, n_5206);
  not g10863 (n_5207, n5897);
  not g10864 (n_5208, n5901);
  and g10865 (n5902, n_5207, n_5208);
  not g10866 (n_5209, n5902);
  and g10867 (n5903, \a[47] , n_5209);
  and g10868 (n5904, \a[3] , n5903);
  and g10869 (n5905, n_5207, n_5209);
  and g10870 (n5906, \a[4] , \a[46] );
  and g10871 (n5907, \a[17] , \a[33] );
  not g10872 (n_5210, n5906);
  not g10873 (n_5211, n5907);
  and g10874 (n5908, n_5210, n_5211);
  not g10875 (n_5212, n5908);
  and g10876 (n5909, n5905, n_5212);
  not g10877 (n_5213, n5904);
  not g10878 (n_5214, n5909);
  and g10879 (n5910, n_5213, n_5214);
  not g10880 (n_5215, n5895);
  not g10881 (n_5216, n5910);
  and g10882 (n5911, n_5215, n_5216);
  not g10883 (n_5217, n5911);
  and g10884 (n5912, n_5215, n_5217);
  and g10885 (n5913, n_5216, n_5217);
  not g10886 (n_5218, n5912);
  not g10887 (n_5219, n5913);
  and g10888 (n5914, n_5218, n_5219);
  and g10889 (n5915, n1494, n2617);
  and g10890 (n5916, n1492, n3452);
  and g10891 (n5917, n1490, n2865);
  not g10892 (n_5220, n5916);
  not g10893 (n_5221, n5917);
  and g10894 (n5918, n_5220, n_5221);
  not g10895 (n_5222, n5915);
  not g10896 (n_5223, n5918);
  and g10897 (n5919, n_5222, n_5223);
  not g10898 (n_5224, n5919);
  and g10899 (n5920, \a[31] , n_5224);
  and g10900 (n5921, \a[19] , n5920);
  and g10901 (n5922, n_5222, n_5224);
  and g10902 (n5923, \a[20] , \a[30] );
  and g10903 (n5924, \a[21] , \a[29] );
  not g10904 (n_5225, n5923);
  not g10905 (n_5226, n5924);
  and g10906 (n5925, n_5225, n_5226);
  not g10907 (n_5227, n5925);
  and g10908 (n5926, n5922, n_5227);
  not g10909 (n_5228, n5921);
  not g10910 (n_5229, n5926);
  and g10911 (n5927, n_5228, n_5229);
  not g10912 (n_5230, n5914);
  not g10913 (n_5231, n5927);
  and g10914 (n5928, n_5230, n_5231);
  not g10915 (n_5232, n5928);
  and g10916 (n5929, n_5230, n_5232);
  and g10917 (n5930, n_5231, n_5232);
  not g10918 (n_5233, n5929);
  not g10919 (n_5234, n5930);
  and g10920 (n5931, n_5233, n_5234);
  and g10921 (n5932, n335, n5296);
  and g10922 (n5933, \a[36] , \a[44] );
  and g10923 (n5934, n1115, n5933);
  not g10924 (n_5235, n5932);
  not g10925 (n_5236, n5934);
  and g10926 (n5935, n_5235, n_5236);
  and g10927 (n5936, \a[7] , \a[43] );
  and g10928 (n5937, \a[14] , \a[36] );
  and g10929 (n5938, n5936, n5937);
  not g10930 (n_5237, n5935);
  not g10931 (n_5238, n5938);
  and g10932 (n5939, n_5237, n_5238);
  not g10933 (n_5239, n5939);
  and g10934 (n5940, n_5238, n_5239);
  not g10935 (n_5240, n5936);
  not g10936 (n_5241, n5937);
  and g10937 (n5941, n_5240, n_5241);
  not g10938 (n_5242, n5941);
  and g10939 (n5942, n5940, n_5242);
  and g10940 (n5943, \a[44] , n_5239);
  and g10941 (n5944, \a[6] , n5943);
  not g10942 (n_5243, n5942);
  not g10943 (n_5244, n5944);
  and g10944 (n5945, n_5243, n_5244);
  and g10945 (n5946, \a[37] , \a[41] );
  and g10946 (n5947, n526, n5946);
  and g10947 (n5948, n432, n5344);
  and g10948 (n5949, \a[13] , \a[42] );
  and g10949 (n5950, n4830, n5949);
  not g10950 (n_5245, n5948);
  not g10951 (n_5246, n5950);
  and g10952 (n5951, n_5245, n_5246);
  not g10953 (n_5247, n5947);
  not g10954 (n_5248, n5951);
  and g10955 (n5952, n_5247, n_5248);
  not g10956 (n_5249, n5952);
  and g10957 (n5953, \a[42] , n_5249);
  and g10958 (n5954, \a[8] , n5953);
  and g10959 (n5955, n_5247, n_5249);
  and g10960 (n5956, \a[9] , \a[41] );
  not g10961 (n_5250, n3689);
  not g10962 (n_5251, n5956);
  and g10963 (n5957, n_5250, n_5251);
  not g10964 (n_5252, n5957);
  and g10965 (n5958, n5955, n_5252);
  not g10966 (n_5253, n5954);
  not g10967 (n_5254, n5958);
  and g10968 (n5959, n_5253, n_5254);
  not g10969 (n_5255, n5945);
  not g10970 (n_5256, n5959);
  and g10971 (n5960, n_5255, n_5256);
  not g10972 (n_5257, n5960);
  and g10973 (n5961, n_5255, n_5257);
  and g10974 (n5962, n_5256, n_5257);
  not g10975 (n_5258, n5961);
  not g10976 (n_5259, n5962);
  and g10977 (n5963, n_5258, n_5259);
  and g10978 (n5964, n723, n4171);
  and g10979 (n5965, n480, n3803);
  and g10980 (n5966, n602, n5083);
  not g10981 (n_5260, n5965);
  not g10982 (n_5261, n5966);
  and g10983 (n5967, n_5260, n_5261);
  not g10984 (n_5262, n5964);
  not g10985 (n_5263, n5967);
  and g10986 (n5968, n_5262, n_5263);
  not g10987 (n_5264, n5968);
  and g10988 (n5969, \a[38] , n_5264);
  and g10989 (n5970, \a[12] , n5969);
  and g10990 (n5971, n_5262, n_5264);
  and g10991 (n5972, \a[10] , \a[40] );
  not g10992 (n_5265, n5315);
  not g10993 (n_5266, n5972);
  and g10994 (n5973, n_5265, n_5266);
  not g10995 (n_5267, n5973);
  and g10996 (n5974, n5971, n_5267);
  not g10997 (n_5268, n5970);
  not g10998 (n_5269, n5974);
  and g10999 (n5975, n_5268, n_5269);
  not g11000 (n_5270, n5963);
  not g11001 (n_5271, n5975);
  and g11002 (n5976, n_5270, n_5271);
  not g11003 (n_5272, n5976);
  and g11004 (n5977, n_5270, n_5272);
  and g11005 (n5978, n_5271, n_5272);
  not g11006 (n_5273, n5977);
  not g11007 (n_5274, n5978);
  and g11008 (n5979, n_5273, n_5274);
  not g11009 (n_5275, n5931);
  and g11010 (n5980, n_5275, n5979);
  not g11011 (n_5276, n5979);
  and g11012 (n5981, n5931, n_5276);
  not g11013 (n_5277, n5980);
  not g11014 (n_5278, n5981);
  and g11015 (n5982, n_5277, n_5278);
  not g11016 (n_5279, n5982);
  and g11017 (n5983, n5884, n_5279);
  not g11018 (n_5280, n5884);
  and g11019 (n5984, n_5280, n5982);
  not g11020 (n_5281, n5983);
  not g11021 (n_5282, n5984);
  and g11022 (n5985, n_5281, n_5282);
  not g11023 (n_5283, n5847);
  and g11024 (n5986, n_5283, n5985);
  not g11025 (n_5284, n5986);
  and g11026 (n5987, n_5283, n_5284);
  and g11027 (n5988, n5985, n_5284);
  not g11028 (n_5285, n5987);
  not g11029 (n_5286, n5988);
  and g11030 (n5989, n_5285, n_5286);
  not g11031 (n_5287, n5846);
  not g11032 (n_5288, n5989);
  and g11033 (n5990, n_5287, n_5288);
  and g11034 (n5991, n5846, n_5286);
  and g11035 (n5992, n_5285, n5991);
  not g11036 (n_5289, n5990);
  not g11037 (n_5290, n5992);
  and g11038 (n5993, n_5289, n_5290);
  not g11039 (n_5291, n5845);
  and g11040 (n5994, n_5291, n5993);
  not g11041 (n_5292, n5993);
  and g11042 (n5995, n5845, n_5292);
  not g11043 (n_5293, n5994);
  not g11044 (n_5294, n5995);
  and g11045 (n5996, n_5293, n_5294);
  and g11046 (n5997, n_5068, n_5072);
  and g11047 (n5998, n_5110, n_5114);
  and g11048 (n5999, n_5140, n_5144);
  and g11049 (n6000, n5998, n5999);
  not g11050 (n_5295, n5998);
  not g11051 (n_5296, n5999);
  and g11052 (n6001, n_5295, n_5296);
  not g11053 (n_5297, n6000);
  not g11054 (n_5298, n6001);
  and g11055 (n6002, n_5297, n_5298);
  and g11056 (n6003, n_5102, n_5106);
  and g11057 (n6004, n_5122, n_5126);
  and g11058 (n6005, n6003, n6004);
  not g11059 (n_5299, n6003);
  not g11060 (n_5300, n6004);
  and g11061 (n6006, n_5299, n_5300);
  not g11062 (n_5301, n6005);
  not g11063 (n_5302, n6006);
  and g11064 (n6007, n_5301, n_5302);
  and g11065 (n6008, n5671, n5719);
  not g11066 (n_5303, n5671);
  not g11067 (n_5304, n5719);
  and g11068 (n6009, n_5303, n_5304);
  not g11069 (n_5305, n6008);
  not g11070 (n_5306, n6009);
  and g11071 (n6010, n_5305, n_5306);
  not g11072 (n_5307, n6010);
  and g11073 (n6011, n5657, n_5307);
  not g11074 (n_5308, n5657);
  and g11075 (n6012, n_5308, n6010);
  not g11076 (n_5309, n6011);
  not g11077 (n_5310, n6012);
  and g11078 (n6013, n_5309, n_5310);
  and g11079 (n6014, n6007, n6013);
  not g11080 (n_5311, n6007);
  not g11081 (n_5312, n6013);
  and g11082 (n6015, n_5311, n_5312);
  not g11083 (n_5313, n6014);
  not g11084 (n_5314, n6015);
  and g11085 (n6016, n_5313, n_5314);
  and g11086 (n6017, n6002, n6016);
  not g11087 (n_5315, n6002);
  not g11088 (n_5316, n6016);
  and g11089 (n6018, n_5315, n_5316);
  not g11090 (n_5317, n6017);
  not g11091 (n_5318, n6018);
  and g11092 (n6019, n_5317, n_5318);
  not g11093 (n_5319, n6019);
  and g11094 (n6020, n5997, n_5319);
  not g11095 (n_5320, n5997);
  and g11096 (n6021, n_5320, n6019);
  not g11097 (n_5321, n6020);
  not g11098 (n_5322, n6021);
  and g11099 (n6022, n_5321, n_5322);
  and g11100 (n6023, n_5011, n_5026);
  and g11101 (n6024, n_5040, n_5041);
  not g11102 (n_5323, n6024);
  and g11103 (n6025, n_5056, n_5323);
  and g11104 (n6026, n6023, n6025);
  not g11105 (n_5324, n6023);
  not g11106 (n_5325, n6025);
  and g11107 (n6027, n_5324, n_5325);
  not g11108 (n_5326, n6026);
  not g11109 (n_5327, n6027);
  and g11110 (n6028, n_5326, n_5327);
  and g11111 (n6029, \a[1] , \a[49] );
  and g11112 (n6030, n2301, n6029);
  not g11113 (n_5328, n2301);
  not g11114 (n_5329, n6029);
  and g11115 (n6031, n_5328, n_5329);
  not g11116 (n_5330, n6030);
  not g11117 (n_5331, n6031);
  and g11118 (n6032, n_5330, n_5331);
  not g11119 (n_5332, n6032);
  and g11120 (n6033, n5638, n_5332);
  not g11121 (n_5333, n5638);
  and g11122 (n6034, n_5333, n6032);
  not g11123 (n_5334, n6033);
  not g11124 (n_5335, n6034);
  and g11125 (n6035, n_5334, n_5335);
  not g11126 (n_5336, n5701);
  and g11127 (n6036, n_5336, n6035);
  not g11128 (n_5337, n6035);
  and g11129 (n6037, n5701, n_5337);
  not g11130 (n_5338, n6036);
  not g11131 (n_5339, n6037);
  and g11132 (n6038, n_5338, n_5339);
  and g11133 (n6039, n6028, n6038);
  not g11134 (n_5340, n6028);
  not g11135 (n_5341, n6038);
  and g11136 (n6040, n_5340, n_5341);
  not g11137 (n_5342, n6039);
  not g11138 (n_5343, n6040);
  and g11139 (n6041, n_5342, n_5343);
  and g11140 (n6042, n5683, n5736);
  not g11141 (n_5344, n5683);
  not g11142 (n_5345, n5736);
  and g11143 (n6043, n_5344, n_5345);
  not g11144 (n_5346, n6042);
  not g11145 (n_5347, n6043);
  and g11146 (n6044, n_5346, n_5347);
  not g11147 (n_5348, n6044);
  and g11148 (n6045, n5626, n_5348);
  not g11149 (n_5349, n5626);
  and g11150 (n6046, n_5349, n6044);
  not g11151 (n_5350, n6045);
  not g11152 (n_5351, n6046);
  and g11153 (n6047, n_5350, n_5351);
  and g11154 (n6048, n_4974, n_4989);
  not g11155 (n_5352, n6047);
  and g11156 (n6049, n_5352, n6048);
  not g11157 (n_5353, n6048);
  and g11158 (n6050, n6047, n_5353);
  not g11159 (n_5354, n6049);
  not g11160 (n_5355, n6050);
  and g11161 (n6051, n_5354, n_5355);
  and g11162 (n6052, n_5081, n_5085);
  not g11163 (n_5356, n6051);
  and g11164 (n6053, n_5356, n6052);
  not g11165 (n_5357, n6052);
  and g11166 (n6054, n6051, n_5357);
  not g11167 (n_5358, n6053);
  not g11168 (n_5359, n6054);
  and g11169 (n6055, n_5358, n_5359);
  and g11170 (n6056, n_5058, n5744);
  not g11171 (n_5360, n6056);
  and g11172 (n6057, n_5064, n_5360);
  not g11173 (n_5361, n6057);
  and g11174 (n6058, n6055, n_5361);
  not g11175 (n_5362, n6055);
  and g11176 (n6059, n_5362, n6057);
  not g11177 (n_5363, n6058);
  not g11178 (n_5364, n6059);
  and g11179 (n6060, n_5363, n_5364);
  and g11180 (n6061, n6041, n6060);
  not g11181 (n_5365, n6041);
  not g11182 (n_5366, n6060);
  and g11183 (n6062, n_5365, n_5366);
  not g11184 (n_5367, n6061);
  not g11185 (n_5368, n6062);
  and g11186 (n6063, n_5367, n_5368);
  and g11187 (n6064, n6022, n6063);
  not g11188 (n_5369, n6022);
  not g11189 (n_5370, n6063);
  and g11190 (n6065, n_5369, n_5370);
  not g11191 (n_5371, n6064);
  not g11192 (n_5372, n6065);
  and g11193 (n6066, n_5371, n_5372);
  and g11194 (n6067, n5996, n6066);
  not g11195 (n_5373, n5996);
  not g11196 (n_5374, n6066);
  and g11197 (n6068, n_5373, n_5374);
  not g11198 (n_5375, n6067);
  not g11199 (n_5376, n6068);
  and g11200 (n6069, n_5375, n_5376);
  not g11201 (n_5377, n6069);
  and g11202 (n6070, n5844, n_5377);
  not g11203 (n_5378, n5844);
  and g11204 (n6071, n_5378, n6069);
  not g11205 (n_5379, n6070);
  not g11206 (n_5380, n6071);
  and g11207 (n6072, n_5379, n_5380);
  not g11208 (n_5381, n6072);
  and g11209 (n6073, n5843, n_5381);
  not g11210 (n_5382, n5843);
  and g11211 (n6074, n_5382, n_5379);
  and g11212 (n6075, n_5380, n6074);
  not g11213 (n_5383, n6073);
  not g11214 (n_5384, n6075);
  and g11215 (\asquared[51] , n_5383, n_5384);
  not g11216 (n_5385, n6074);
  and g11217 (n6077, n_5380, n_5385);
  and g11218 (n6078, n_5293, n_5375);
  and g11219 (n6079, n_5322, n_5371);
  and g11220 (n6080, n_5363, n_5367);
  and g11221 (n6081, n_5298, n_5317);
  and g11222 (n6082, \a[0] , \a[51] );
  and g11223 (n6083, n6030, n6082);
  not g11224 (n_5387, n6083);
  and g11225 (n6084, n6030, n_5387);
  and g11226 (n6085, n_5330, n6082);
  not g11227 (n_5388, n6084);
  not g11228 (n_5389, n6085);
  and g11229 (n6086, n_5388, n_5389);
  and g11230 (n6087, \a[1] , \a[50] );
  and g11231 (n6088, \a[26] , n6087);
  not g11232 (n_5390, n6088);
  and g11233 (n6089, \a[26] , n_5390);
  and g11234 (n6090, n6087, n_5390);
  not g11235 (n_5391, n6089);
  not g11236 (n_5392, n6090);
  and g11237 (n6091, n_5391, n_5392);
  not g11238 (n_5393, n6086);
  not g11239 (n_5394, n6091);
  and g11240 (n6092, n_5393, n_5394);
  not g11241 (n_5395, n6092);
  and g11242 (n6093, n_5393, n_5395);
  and g11243 (n6094, n_5394, n_5395);
  not g11244 (n_5396, n6093);
  not g11245 (n_5397, n6094);
  and g11246 (n6095, n_5396, n_5397);
  and g11247 (n6096, n1490, n3812);
  not g11248 (n_5398, n6096);
  and g11250 (n6098, \a[20] , \a[31] );
  and g11251 (n6099, \a[19] , \a[32] );
  not g11252 (n_5399, n6098);
  not g11253 (n_5400, n6099);
  and g11254 (n6100, n_5399, n_5400);
  not g11255 (n_5401, n6100);
  not g11258 (n_5402, n6102);
  and g11259 (n6103, \a[34] , n_5402);
  and g11260 (n6104, \a[17] , n6103);
  and g11261 (n6105, n_5398, n_5402);
  and g11262 (n6106, n_5401, n6105);
  not g11263 (n_5403, n6104);
  not g11264 (n_5404, n6106);
  and g11265 (n6107, n_5403, n_5404);
  not g11266 (n_5405, n6095);
  not g11267 (n_5406, n6107);
  and g11268 (n6108, n_5405, n_5406);
  not g11269 (n_5407, n6108);
  and g11270 (n6109, n_5405, n_5407);
  and g11271 (n6110, n_5406, n_5407);
  not g11272 (n_5408, n6109);
  not g11273 (n_5409, n6110);
  and g11274 (n6111, n_5408, n_5409);
  and g11275 (n6112, n_5347, n_5351);
  and g11276 (n6113, n6111, n6112);
  not g11277 (n_5410, n6111);
  not g11278 (n_5411, n6112);
  and g11279 (n6114, n_5410, n_5411);
  not g11280 (n_5412, n6113);
  not g11281 (n_5413, n6114);
  and g11282 (n6115, n_5412, n_5413);
  and g11283 (n6116, n1340, n5896);
  and g11284 (n6117, n1050, n2972);
  not g11285 (n_5414, n6116);
  not g11286 (n_5415, n6117);
  and g11287 (n6118, n_5414, n_5415);
  and g11288 (n6119, \a[5] , \a[46] );
  and g11289 (n6120, \a[16] , \a[35] );
  and g11290 (n6121, n6119, n6120);
  not g11291 (n_5416, n6118);
  not g11292 (n_5417, n6121);
  and g11293 (n6122, n_5416, n_5417);
  not g11294 (n_5418, n6122);
  and g11295 (n6123, n_5417, n_5418);
  not g11296 (n_5419, n6119);
  not g11297 (n_5420, n6120);
  and g11298 (n6124, n_5419, n_5420);
  not g11299 (n_5421, n6124);
  and g11300 (n6125, n6123, n_5421);
  and g11301 (n6126, \a[33] , n_5418);
  and g11302 (n6127, \a[18] , n6126);
  not g11303 (n_5422, n6125);
  not g11304 (n_5423, n6127);
  and g11305 (n6128, n_5422, n_5423);
  and g11306 (n6129, n1919, n2334);
  and g11307 (n6130, n1367, n3110);
  and g11308 (n6131, n1574, n2617);
  not g11309 (n_5424, n6130);
  not g11310 (n_5425, n6131);
  and g11311 (n6132, n_5424, n_5425);
  not g11312 (n_5426, n6129);
  not g11313 (n_5427, n6132);
  and g11314 (n6133, n_5426, n_5427);
  not g11315 (n_5428, n6133);
  and g11316 (n6134, \a[30] , n_5428);
  and g11317 (n6135, \a[21] , n6134);
  and g11318 (n6136, \a[22] , \a[29] );
  and g11319 (n6137, \a[23] , \a[28] );
  not g11320 (n_5429, n6136);
  not g11321 (n_5430, n6137);
  and g11322 (n6138, n_5429, n_5430);
  and g11323 (n6139, n_5426, n_5428);
  not g11324 (n_5431, n6138);
  and g11325 (n6140, n_5431, n6139);
  not g11326 (n_5432, n6135);
  not g11327 (n_5433, n6140);
  and g11328 (n6141, n_5432, n_5433);
  not g11329 (n_5434, n6128);
  not g11330 (n_5435, n6141);
  and g11331 (n6142, n_5434, n_5435);
  not g11332 (n_5436, n6142);
  and g11333 (n6143, n_5434, n_5436);
  and g11334 (n6144, n_5435, n_5436);
  not g11335 (n_5437, n6143);
  not g11336 (n_5438, n6144);
  and g11337 (n6145, n_5437, n_5438);
  and g11338 (n6146, \a[37] , \a[45] );
  and g11339 (n6147, n1115, n6146);
  and g11340 (n6148, \a[6] , \a[45] );
  and g11341 (n6149, \a[36] , n6148);
  and g11342 (n6150, \a[15] , n6149);
  and g11343 (n6151, n895, n3687);
  not g11344 (n_5439, n6150);
  not g11345 (n_5440, n6151);
  and g11346 (n6152, n_5439, n_5440);
  not g11347 (n_5441, n6147);
  not g11348 (n_5442, n6152);
  and g11349 (n6153, n_5441, n_5442);
  not g11350 (n_5443, n6153);
  and g11351 (n6154, \a[36] , n_5443);
  and g11352 (n6155, \a[15] , n6154);
  and g11353 (n6156, \a[14] , \a[37] );
  not g11354 (n_5444, n6148);
  not g11355 (n_5445, n6156);
  and g11356 (n6157, n_5444, n_5445);
  and g11357 (n6158, n_5441, n_5443);
  not g11358 (n_5446, n6157);
  and g11359 (n6159, n_5446, n6158);
  not g11360 (n_5447, n6155);
  not g11361 (n_5448, n6159);
  and g11362 (n6160, n_5447, n_5448);
  not g11363 (n_5449, n6145);
  not g11364 (n_5450, n6160);
  and g11365 (n6161, n_5449, n_5450);
  not g11366 (n_5451, n6161);
  and g11367 (n6162, n_5449, n_5451);
  and g11368 (n6163, n_5450, n_5451);
  not g11369 (n_5452, n6162);
  not g11370 (n_5453, n6163);
  and g11371 (n6164, n_5452, n_5453);
  and g11372 (n6165, \a[13] , \a[43] );
  and g11373 (n6166, n5081, n6165);
  and g11374 (n6167, n380, n5296);
  and g11375 (n6168, \a[13] , \a[44] );
  and g11376 (n6169, n4823, n6168);
  not g11377 (n_5454, n6167);
  not g11378 (n_5455, n6169);
  and g11379 (n6170, n_5454, n_5455);
  not g11380 (n_5456, n6166);
  not g11381 (n_5457, n6170);
  and g11382 (n6171, n_5456, n_5457);
  not g11383 (n_5458, n6171);
  and g11384 (n6172, n_5456, n_5458);
  and g11385 (n6173, \a[8] , \a[43] );
  and g11386 (n6174, \a[13] , \a[38] );
  not g11387 (n_5459, n6173);
  not g11388 (n_5460, n6174);
  and g11389 (n6175, n_5459, n_5460);
  not g11390 (n_5461, n6175);
  and g11391 (n6176, n6172, n_5461);
  and g11392 (n6177, \a[44] , n_5458);
  and g11393 (n6178, \a[7] , n6177);
  not g11394 (n_5462, n6176);
  not g11395 (n_5463, n6178);
  and g11396 (n6179, n_5462, n_5463);
  and g11397 (n6180, \a[9] , \a[42] );
  and g11398 (n6181, n480, n3984);
  and g11399 (n6182, n4750, n6180);
  and g11400 (n6183, n484, n5344);
  not g11401 (n_5464, n6182);
  not g11402 (n_5465, n6183);
  and g11403 (n6184, n_5464, n_5465);
  not g11404 (n_5466, n6181);
  not g11405 (n_5467, n6184);
  and g11406 (n6185, n_5466, n_5467);
  not g11407 (n_5468, n6185);
  and g11408 (n6186, n6180, n_5468);
  and g11409 (n6187, n_5466, n_5468);
  and g11410 (n6188, \a[10] , \a[41] );
  not g11411 (n_5469, n4750);
  not g11412 (n_5470, n6188);
  and g11413 (n6189, n_5469, n_5470);
  not g11414 (n_5471, n6189);
  and g11415 (n6190, n6187, n_5471);
  not g11416 (n_5472, n6186);
  not g11417 (n_5473, n6190);
  and g11418 (n6191, n_5472, n_5473);
  not g11419 (n_5474, n6179);
  not g11420 (n_5475, n6191);
  and g11421 (n6192, n_5474, n_5475);
  not g11422 (n_5476, n6192);
  and g11423 (n6193, n_5474, n_5476);
  and g11424 (n6194, n_5475, n_5476);
  not g11425 (n_5477, n6193);
  not g11426 (n_5478, n6194);
  and g11427 (n6195, n_5477, n_5478);
  and g11428 (n6196, \a[24] , \a[27] );
  not g11429 (n_5479, n2463);
  not g11430 (n_5480, n6196);
  and g11431 (n6197, n_5479, n_5480);
  and g11432 (n6198, n1904, n2227);
  not g11433 (n_5481, n6198);
  not g11436 (n_5482, n6197);
  not g11438 (n_5483, n6201);
  and g11439 (n6202, \a[40] , n_5483);
  and g11440 (n6203, \a[11] , n6202);
  and g11441 (n6204, n_5481, n_5483);
  and g11442 (n6205, n_5482, n6204);
  not g11443 (n_5484, n6203);
  not g11444 (n_5485, n6205);
  and g11445 (n6206, n_5484, n_5485);
  not g11446 (n_5486, n6195);
  not g11447 (n_5487, n6206);
  and g11448 (n6207, n_5486, n_5487);
  not g11449 (n_5488, n6207);
  and g11450 (n6208, n_5486, n_5488);
  and g11451 (n6209, n_5487, n_5488);
  not g11452 (n_5489, n6208);
  not g11453 (n_5490, n6209);
  and g11454 (n6210, n_5489, n_5490);
  not g11455 (n_5491, n6164);
  and g11456 (n6211, n_5491, n6210);
  not g11457 (n_5492, n6210);
  and g11458 (n6212, n6164, n_5492);
  not g11459 (n_5493, n6211);
  not g11460 (n_5494, n6212);
  and g11461 (n6213, n_5493, n_5494);
  not g11462 (n_5495, n6213);
  and g11463 (n6214, n6115, n_5495);
  not g11464 (n_5496, n6115);
  and g11465 (n6215, n_5496, n6213);
  not g11466 (n_5497, n6214);
  not g11467 (n_5498, n6215);
  and g11468 (n6216, n_5497, n_5498);
  not g11469 (n_5499, n6081);
  and g11470 (n6217, n_5499, n6216);
  not g11471 (n_5500, n6216);
  and g11472 (n6218, n6081, n_5500);
  not g11473 (n_5501, n6217);
  not g11474 (n_5502, n6218);
  and g11475 (n6219, n_5501, n_5502);
  not g11476 (n_5503, n6080);
  and g11477 (n6220, n_5503, n6219);
  not g11478 (n_5504, n6219);
  and g11479 (n6221, n6080, n_5504);
  not g11480 (n_5505, n6220);
  not g11481 (n_5506, n6221);
  and g11482 (n6222, n_5505, n_5506);
  not g11483 (n_5507, n6079);
  and g11484 (n6223, n_5507, n6222);
  not g11485 (n_5508, n6222);
  and g11486 (n6224, n6079, n_5508);
  not g11487 (n_5509, n6223);
  not g11488 (n_5510, n6224);
  and g11489 (n6225, n_5509, n_5510);
  and g11490 (n6226, n_5284, n_5289);
  and g11491 (n6227, n_5355, n_5359);
  and g11492 (n6228, n_5327, n_5342);
  and g11493 (n6229, n6227, n6228);
  not g11494 (n_5511, n6227);
  not g11495 (n_5512, n6228);
  and g11496 (n6230, n_5511, n_5512);
  not g11497 (n_5513, n6229);
  not g11498 (n_5514, n6230);
  and g11499 (n6231, n_5513, n_5514);
  and g11500 (n6232, n_5306, n_5310);
  and g11501 (n6233, n_5335, n_5338);
  and g11502 (n6234, n6232, n6233);
  not g11503 (n_5515, n6232);
  not g11504 (n_5516, n6233);
  and g11505 (n6235, n_5515, n_5516);
  not g11506 (n_5517, n6234);
  not g11507 (n_5518, n6235);
  and g11508 (n6236, n_5517, n_5518);
  and g11509 (n6237, n_5217, n_5232);
  not g11510 (n_5519, n6236);
  and g11511 (n6238, n_5519, n6237);
  not g11512 (n_5520, n6237);
  and g11513 (n6239, n6236, n_5520);
  not g11514 (n_5521, n6238);
  not g11515 (n_5522, n6239);
  and g11516 (n6240, n_5521, n_5522);
  and g11517 (n6241, n6231, n6240);
  not g11518 (n_5523, n6231);
  not g11519 (n_5524, n6240);
  and g11520 (n6242, n_5523, n_5524);
  not g11521 (n_5525, n6241);
  not g11522 (n_5526, n6242);
  and g11523 (n6243, n_5525, n_5526);
  not g11524 (n_5527, n6226);
  and g11525 (n6244, n_5527, n6243);
  not g11526 (n_5528, n6243);
  and g11527 (n6245, n6226, n_5528);
  not g11528 (n_5529, n6244);
  not g11529 (n_5530, n6245);
  and g11530 (n6246, n_5529, n_5530);
  and g11531 (n6247, n_5275, n_5276);
  not g11532 (n_5531, n6247);
  and g11533 (n6248, n_5281, n_5531);
  and g11534 (n6249, n5855, n5971);
  not g11535 (n_5532, n5855);
  not g11536 (n_5533, n5971);
  and g11537 (n6250, n_5532, n_5533);
  not g11538 (n_5534, n6249);
  not g11539 (n_5535, n6250);
  and g11540 (n6251, n_5534, n_5535);
  and g11541 (n6252, \a[47] , \a[48] );
  and g11542 (n6253, n209, n6252);
  and g11543 (n6254, \a[47] , \a[49] );
  and g11544 (n6255, n252, n6254);
  and g11545 (n6256, \a[48] , \a[49] );
  and g11546 (n6257, n218, n6256);
  not g11547 (n_5536, n6255);
  not g11548 (n_5537, n6257);
  and g11549 (n6258, n_5536, n_5537);
  not g11550 (n_5538, n6253);
  not g11551 (n_5539, n6258);
  and g11552 (n6259, n_5538, n_5539);
  not g11553 (n_5540, n6259);
  and g11554 (n6260, \a[49] , n_5540);
  and g11555 (n6261, \a[2] , n6260);
  and g11556 (n6262, n_5538, n_5540);
  and g11557 (n6263, \a[3] , \a[48] );
  and g11558 (n6264, \a[4] , \a[47] );
  not g11559 (n_5541, n6263);
  not g11560 (n_5542, n6264);
  and g11561 (n6265, n_5541, n_5542);
  not g11562 (n_5543, n6265);
  and g11563 (n6266, n6262, n_5543);
  not g11564 (n_5544, n6261);
  not g11565 (n_5545, n6266);
  and g11566 (n6267, n_5544, n_5545);
  not g11567 (n_5546, n6267);
  and g11568 (n6268, n6251, n_5546);
  not g11569 (n_5547, n6268);
  and g11570 (n6269, n6251, n_5547);
  and g11571 (n6270, n_5546, n_5547);
  not g11572 (n_5548, n6269);
  not g11573 (n_5549, n6270);
  and g11574 (n6271, n_5548, n_5549);
  and g11575 (n6272, n_5190, n_5196);
  and g11576 (n6273, n6271, n6272);
  not g11577 (n_5550, n6271);
  not g11578 (n_5551, n6272);
  and g11579 (n6274, n_5550, n_5551);
  not g11580 (n_5552, n6273);
  not g11581 (n_5553, n6274);
  and g11582 (n6275, n_5552, n_5553);
  and g11583 (n6276, n_5302, n_5313);
  not g11584 (n_5554, n6276);
  and g11585 (n6277, n6275, n_5554);
  not g11586 (n_5555, n6275);
  and g11587 (n6278, n_5555, n6276);
  not g11588 (n_5556, n6277);
  not g11589 (n_5557, n6278);
  and g11590 (n6279, n_5556, n_5557);
  not g11591 (n_5558, n6248);
  and g11592 (n6280, n_5558, n6279);
  not g11593 (n_5559, n6279);
  and g11594 (n6281, n6248, n_5559);
  not g11595 (n_5560, n6280);
  not g11596 (n_5561, n6281);
  and g11597 (n6282, n_5560, n_5561);
  and g11598 (n6283, n5940, n5955);
  not g11599 (n_5562, n5940);
  not g11600 (n_5563, n5955);
  and g11601 (n6284, n_5562, n_5563);
  not g11602 (n_5564, n6283);
  not g11603 (n_5565, n6284);
  and g11604 (n6285, n_5564, n_5565);
  not g11605 (n_5566, n6285);
  and g11606 (n6286, n5874, n_5566);
  not g11607 (n_5567, n5874);
  and g11608 (n6287, n_5567, n6285);
  not g11609 (n_5568, n6286);
  not g11610 (n_5569, n6287);
  and g11611 (n6288, n_5568, n_5569);
  and g11612 (n6289, n_5257, n_5272);
  not g11613 (n_5570, n6288);
  and g11614 (n6290, n_5570, n6289);
  not g11615 (n_5571, n6289);
  and g11616 (n6291, n6288, n_5571);
  not g11617 (n_5572, n6290);
  not g11618 (n_5573, n6291);
  and g11619 (n6292, n_5572, n_5573);
  and g11620 (n6293, n5905, n5922);
  not g11621 (n_5574, n5905);
  not g11622 (n_5575, n5922);
  and g11623 (n6294, n_5574, n_5575);
  not g11624 (n_5576, n6293);
  not g11625 (n_5577, n6294);
  and g11626 (n6295, n_5576, n_5577);
  not g11627 (n_5578, n6295);
  and g11628 (n6296, n5892, n_5578);
  not g11629 (n_5579, n5892);
  and g11630 (n6297, n_5579, n6295);
  not g11631 (n_5580, n6296);
  not g11632 (n_5581, n6297);
  and g11633 (n6298, n_5580, n_5581);
  and g11634 (n6299, n6292, n6298);
  not g11635 (n_5582, n6292);
  not g11636 (n_5583, n6298);
  and g11637 (n6300, n_5582, n_5583);
  not g11638 (n_5584, n6299);
  not g11639 (n_5585, n6300);
  and g11640 (n6301, n_5584, n_5585);
  and g11641 (n6302, n6282, n6301);
  not g11642 (n_5586, n6282);
  not g11643 (n_5587, n6301);
  and g11644 (n6303, n_5586, n_5587);
  not g11645 (n_5588, n6302);
  not g11646 (n_5589, n6303);
  and g11647 (n6304, n_5588, n_5589);
  and g11648 (n6305, n6246, n6304);
  not g11649 (n_5590, n6246);
  not g11650 (n_5591, n6304);
  and g11651 (n6306, n_5590, n_5591);
  not g11652 (n_5592, n6305);
  not g11653 (n_5593, n6306);
  and g11654 (n6307, n_5592, n_5593);
  and g11655 (n6308, n6225, n6307);
  not g11656 (n_5594, n6225);
  not g11657 (n_5595, n6307);
  and g11658 (n6309, n_5594, n_5595);
  not g11659 (n_5596, n6308);
  not g11660 (n_5597, n6309);
  and g11661 (n6310, n_5596, n_5597);
  not g11662 (n_5598, n6078);
  and g11663 (n6311, n_5598, n6310);
  not g11664 (n_5599, n6310);
  and g11665 (n6312, n6078, n_5599);
  not g11666 (n_5600, n6311);
  not g11667 (n_5601, n6312);
  and g11668 (n6313, n_5600, n_5601);
  not g11669 (n_5602, n6077);
  not g11670 (n_5603, n6313);
  and g11671 (n6314, n_5602, n_5603);
  and g11672 (n6315, n6077, n6313);
  or g11673 (\asquared[52] , n6314, n6315);
  and g11674 (n6317, n_5602, n_5601);
  not g11675 (n_5604, n6317);
  and g11676 (n6318, n_5600, n_5604);
  and g11677 (n6319, n_5509, n_5596);
  and g11678 (n6320, n_5501, n_5505);
  and g11679 (n6321, n_5577, n_5581);
  and g11680 (n6322, \a[2] , \a[50] );
  and g11681 (n6323, \a[3] , \a[49] );
  not g11682 (n_5605, n6322);
  not g11683 (n_5606, n6323);
  and g11684 (n6324, n_5605, n_5606);
  and g11685 (n6325, \a[49] , \a[50] );
  and g11686 (n6326, n218, n6325);
  not g11687 (n_5607, n6326);
  not g11690 (n_5608, n6324);
  not g11692 (n_5609, n6329);
  and g11693 (n6330, \a[33] , n_5609);
  and g11694 (n6331, \a[19] , n6330);
  and g11695 (n6332, n_5607, n_5609);
  and g11696 (n6333, n_5608, n6332);
  not g11697 (n_5610, n6331);
  not g11698 (n_5611, n6333);
  and g11699 (n6334, n_5610, n_5611);
  not g11700 (n_5612, n6321);
  not g11701 (n_5613, n6334);
  and g11702 (n6335, n_5612, n_5613);
  not g11703 (n_5614, n6335);
  and g11704 (n6336, n_5612, n_5614);
  and g11705 (n6337, n_5613, n_5614);
  not g11706 (n_5615, n6336);
  not g11707 (n_5616, n6337);
  and g11708 (n6338, n_5615, n_5616);
  and g11709 (n6339, n_5565, n_5569);
  and g11710 (n6340, n6338, n6339);
  not g11711 (n_5617, n6338);
  not g11712 (n_5618, n6339);
  and g11713 (n6341, n_5617, n_5618);
  not g11714 (n_5619, n6340);
  not g11715 (n_5620, n6341);
  and g11716 (n6342, n_5619, n_5620);
  and g11717 (n6343, n_5553, n_5556);
  not g11718 (n_5621, n6342);
  and g11719 (n6344, n_5621, n6343);
  not g11720 (n_5622, n6343);
  and g11721 (n6345, n6342, n_5622);
  not g11722 (n_5623, n6344);
  not g11723 (n_5624, n6345);
  and g11724 (n6346, n_5623, n_5624);
  and g11725 (n6347, n_5476, n_5488);
  and g11726 (n6348, n_5535, n_5547);
  and g11727 (n6349, \a[1] , \a[51] );
  not g11728 (n_5625, n2633);
  not g11729 (n_5626, n6349);
  and g11730 (n6350, n_5625, n_5626);
  and g11731 (n6351, n2633, n6349);
  not g11732 (n_5627, n6350);
  not g11733 (n_5628, n6351);
  and g11734 (n6352, n_5627, n_5628);
  and g11735 (n6353, n6088, n6352);
  not g11736 (n_5629, n6352);
  and g11737 (n6354, n_5390, n_5629);
  not g11738 (n_5630, n6353);
  not g11739 (n_5631, n6354);
  and g11740 (n6355, n_5630, n_5631);
  not g11741 (n_5632, n6204);
  and g11742 (n6356, n_5632, n6355);
  not g11743 (n_5633, n6355);
  and g11744 (n6357, n6204, n_5633);
  not g11745 (n_5634, n6356);
  not g11746 (n_5635, n6357);
  and g11747 (n6358, n_5634, n_5635);
  not g11748 (n_5636, n6348);
  and g11749 (n6359, n_5636, n6358);
  not g11750 (n_5637, n6358);
  and g11751 (n6360, n6348, n_5637);
  not g11752 (n_5638, n6359);
  not g11753 (n_5639, n6360);
  and g11754 (n6361, n_5638, n_5639);
  not g11755 (n_5640, n6347);
  and g11756 (n6362, n_5640, n6361);
  not g11757 (n_5641, n6361);
  and g11758 (n6363, n6347, n_5641);
  not g11759 (n_5642, n6362);
  not g11760 (n_5643, n6363);
  and g11761 (n6364, n_5642, n_5643);
  and g11762 (n6365, n6346, n6364);
  not g11763 (n_5644, n6346);
  not g11764 (n_5645, n6364);
  and g11765 (n6366, n_5644, n_5645);
  not g11766 (n_5646, n6365);
  not g11767 (n_5647, n6366);
  and g11768 (n6367, n_5646, n_5647);
  not g11769 (n_5648, n6367);
  and g11770 (n6368, n6320, n_5648);
  not g11771 (n_5649, n6320);
  and g11772 (n6369, n_5649, n6367);
  not g11773 (n_5650, n6368);
  not g11774 (n_5651, n6369);
  and g11775 (n6370, n_5650, n_5651);
  and g11776 (n6371, n_5387, n_5395);
  and g11777 (n6372, n6187, n6371);
  not g11778 (n_5652, n6187);
  not g11779 (n_5653, n6371);
  and g11780 (n6373, n_5652, n_5653);
  not g11781 (n_5654, n6372);
  not g11782 (n_5655, n6373);
  and g11783 (n6374, n_5654, n_5655);
  and g11784 (n6375, \a[35] , n793);
  and g11785 (n6376, \a[48] , n212);
  not g11786 (n_5656, n6375);
  not g11787 (n_5657, n6376);
  and g11788 (n6377, n_5656, n_5657);
  and g11789 (n6378, \a[4] , \a[48] );
  and g11790 (n6379, \a[17] , \a[35] );
  and g11791 (n6380, n6378, n6379);
  not g11792 (n_5659, n6380);
  and g11793 (n6381, \a[52] , n_5659);
  not g11794 (n_5660, n6377);
  and g11795 (n6382, n_5660, n6381);
  not g11796 (n_5661, n6382);
  and g11797 (n6383, \a[52] , n_5661);
  and g11798 (n6384, \a[0] , n6383);
  and g11799 (n6385, n_5659, n_5661);
  not g11800 (n_5662, n6378);
  not g11801 (n_5663, n6379);
  and g11802 (n6386, n_5662, n_5663);
  not g11803 (n_5664, n6386);
  and g11804 (n6387, n6385, n_5664);
  not g11805 (n_5665, n6384);
  not g11806 (n_5666, n6387);
  and g11807 (n6388, n_5665, n_5666);
  not g11808 (n_5667, n6388);
  and g11809 (n6389, n6374, n_5667);
  not g11810 (n_5668, n6389);
  and g11811 (n6390, n6374, n_5668);
  and g11812 (n6391, n_5667, n_5668);
  not g11813 (n_5669, n6390);
  not g11814 (n_5670, n6391);
  and g11815 (n6392, n_5669, n_5670);
  and g11816 (n6393, n_5407, n_5413);
  and g11817 (n6394, n6392, n6393);
  not g11818 (n_5671, n6392);
  not g11819 (n_5672, n6393);
  and g11820 (n6395, n_5671, n_5672);
  not g11821 (n_5673, n6394);
  not g11822 (n_5674, n6395);
  and g11823 (n6396, n_5673, n_5674);
  and g11824 (n6397, n_5518, n_5522);
  not g11825 (n_5675, n6396);
  and g11826 (n6398, n_5675, n6397);
  not g11827 (n_5676, n6397);
  and g11828 (n6399, n6396, n_5676);
  not g11829 (n_5677, n6398);
  not g11830 (n_5678, n6399);
  and g11831 (n6400, n_5677, n_5678);
  and g11832 (n6401, n_5491, n_5492);
  not g11833 (n_5679, n6401);
  and g11834 (n6402, n_5497, n_5679);
  and g11835 (n6403, n6123, n6172);
  not g11836 (n_5680, n6123);
  not g11837 (n_5681, n6172);
  and g11838 (n6404, n_5680, n_5681);
  not g11839 (n_5682, n6403);
  not g11840 (n_5683, n6404);
  and g11841 (n6405, n_5682, n_5683);
  not g11842 (n_5684, n6405);
  and g11843 (n6406, n6139, n_5684);
  not g11844 (n_5685, n6139);
  and g11845 (n6407, n_5685, n6405);
  not g11846 (n_5686, n6406);
  not g11847 (n_5687, n6407);
  and g11848 (n6408, n_5686, n_5687);
  and g11849 (n6409, n6105, n6262);
  not g11850 (n_5688, n6105);
  not g11851 (n_5689, n6262);
  and g11852 (n6410, n_5688, n_5689);
  not g11853 (n_5690, n6409);
  not g11854 (n_5691, n6410);
  and g11855 (n6411, n_5690, n_5691);
  not g11856 (n_5692, n6411);
  and g11857 (n6412, n6158, n_5692);
  not g11858 (n_5693, n6158);
  and g11859 (n6413, n_5693, n6411);
  not g11860 (n_5694, n6412);
  not g11861 (n_5695, n6413);
  and g11862 (n6414, n_5694, n_5695);
  and g11863 (n6415, n_5436, n_5451);
  not g11864 (n_5696, n6414);
  and g11865 (n6416, n_5696, n6415);
  not g11866 (n_5697, n6415);
  and g11867 (n6417, n6414, n_5697);
  not g11868 (n_5698, n6416);
  not g11869 (n_5699, n6417);
  and g11870 (n6418, n_5698, n_5699);
  and g11871 (n6419, n6408, n6418);
  not g11872 (n_5700, n6408);
  not g11873 (n_5701, n6418);
  and g11874 (n6420, n_5700, n_5701);
  not g11875 (n_5702, n6419);
  not g11876 (n_5703, n6420);
  and g11877 (n6421, n_5702, n_5703);
  not g11878 (n_5704, n6402);
  and g11879 (n6422, n_5704, n6421);
  not g11880 (n_5705, n6422);
  and g11881 (n6423, n_5704, n_5705);
  and g11882 (n6424, n6421, n_5705);
  not g11883 (n_5706, n6423);
  not g11884 (n_5707, n6424);
  and g11885 (n6425, n_5706, n_5707);
  not g11886 (n_5708, n6425);
  and g11887 (n6426, n6400, n_5708);
  not g11888 (n_5709, n6426);
  and g11889 (n6427, n6400, n_5709);
  and g11890 (n6428, n_5708, n_5709);
  not g11891 (n_5710, n6427);
  not g11892 (n_5711, n6428);
  and g11893 (n6429, n_5710, n_5711);
  not g11894 (n_5712, n6429);
  and g11895 (n6430, n6370, n_5712);
  not g11896 (n_5713, n6430);
  and g11897 (n6431, n6370, n_5713);
  and g11898 (n6432, n_5712, n_5713);
  not g11899 (n_5714, n6431);
  not g11900 (n_5715, n6432);
  and g11901 (n6433, n_5714, n_5715);
  and g11902 (n6434, n_5560, n_5588);
  and g11903 (n6435, n_5514, n_5525);
  and g11904 (n6436, n_5573, n_5584);
  and g11905 (n6437, \a[36] , \a[46] );
  and g11906 (n6438, n721, n6437);
  and g11907 (n6439, n332, n5666);
  and g11908 (n6440, \a[5] , \a[47] );
  and g11909 (n6441, \a[16] , \a[36] );
  and g11910 (n6442, n6440, n6441);
  not g11911 (n_5716, n6439);
  not g11912 (n_5717, n6442);
  and g11913 (n6443, n_5716, n_5717);
  not g11914 (n_5718, n6438);
  not g11915 (n_5719, n6443);
  and g11916 (n6444, n_5718, n_5719);
  not g11917 (n_5720, n6444);
  and g11918 (n6445, n_5718, n_5720);
  and g11919 (n6446, \a[6] , \a[46] );
  not g11920 (n_5721, n6441);
  not g11921 (n_5722, n6446);
  and g11922 (n6447, n_5721, n_5722);
  not g11923 (n_5723, n6447);
  and g11924 (n6448, n6445, n_5723);
  and g11925 (n6449, n6440, n_5720);
  not g11926 (n_5724, n6448);
  not g11927 (n_5725, n6449);
  and g11928 (n6450, n_5724, n_5725);
  and g11929 (n6451, \a[10] , \a[42] );
  and g11930 (n6452, n602, n5413);
  and g11931 (n6453, \a[40] , \a[42] );
  and g11932 (n6454, n480, n6453);
  and g11933 (n6455, n723, n5344);
  not g11934 (n_5726, n6454);
  not g11935 (n_5727, n6455);
  and g11936 (n6456, n_5726, n_5727);
  not g11937 (n_5728, n6452);
  not g11938 (n_5729, n6456);
  and g11939 (n6457, n_5728, n_5729);
  not g11940 (n_5730, n6457);
  and g11941 (n6458, n6451, n_5730);
  and g11942 (n6459, n_5728, n_5730);
  and g11943 (n6460, \a[11] , \a[41] );
  not g11944 (n_5731, n5192);
  not g11945 (n_5732, n6460);
  and g11946 (n6461, n_5731, n_5732);
  not g11947 (n_5733, n6461);
  and g11948 (n6462, n6459, n_5733);
  not g11949 (n_5734, n6458);
  not g11950 (n_5735, n6462);
  and g11951 (n6463, n_5734, n_5735);
  not g11952 (n_5736, n6450);
  not g11953 (n_5737, n6463);
  and g11954 (n6464, n_5736, n_5737);
  not g11955 (n_5738, n6464);
  and g11956 (n6465, n_5736, n_5738);
  and g11957 (n6466, n_5737, n_5738);
  not g11958 (n_5739, n6465);
  not g11959 (n_5740, n6466);
  and g11960 (n6467, n_5739, n_5740);
  and g11961 (n6468, \a[7] , \a[45] );
  and g11962 (n6469, \a[8] , \a[44] );
  not g11963 (n_5741, n6468);
  not g11964 (n_5742, n6469);
  and g11965 (n6470, n_5741, n_5742);
  and g11966 (n6471, n380, n5713);
  not g11967 (n_5743, n6471);
  not g11970 (n_5744, n6470);
  not g11972 (n_5745, n6474);
  and g11973 (n6475, \a[37] , n_5745);
  and g11974 (n6476, \a[15] , n6475);
  and g11975 (n6477, n_5743, n_5745);
  and g11976 (n6478, n_5744, n6477);
  not g11977 (n_5746, n6476);
  not g11978 (n_5747, n6478);
  and g11979 (n6479, n_5746, n_5747);
  not g11980 (n_5748, n6467);
  not g11981 (n_5749, n6479);
  and g11982 (n6480, n_5748, n_5749);
  not g11983 (n_5750, n6480);
  and g11984 (n6481, n_5748, n_5750);
  and g11985 (n6482, n_5749, n_5750);
  not g11986 (n_5751, n6481);
  not g11987 (n_5752, n6482);
  and g11988 (n6483, n_5751, n_5752);
  and g11989 (n6484, n1494, n3812);
  and g11990 (n6485, \a[31] , \a[34] );
  and g11991 (n6486, n3648, n6485);
  and g11992 (n6487, n1331, n4090);
  not g11993 (n_5753, n6486);
  not g11994 (n_5754, n6487);
  and g11995 (n6488, n_5753, n_5754);
  not g11996 (n_5755, n6484);
  not g11997 (n_5756, n6488);
  and g11998 (n6489, n_5755, n_5756);
  not g11999 (n_5757, n6489);
  and g12000 (n6490, n_5755, n_5757);
  and g12001 (n6491, \a[20] , \a[32] );
  and g12002 (n6492, \a[21] , \a[31] );
  not g12003 (n_5758, n6491);
  not g12004 (n_5759, n6492);
  and g12005 (n6493, n_5758, n_5759);
  not g12006 (n_5760, n6493);
  and g12007 (n6494, n6490, n_5760);
  and g12008 (n6495, \a[34] , n_5757);
  and g12009 (n6496, \a[18] , n6495);
  not g12010 (n_5761, n6494);
  not g12011 (n_5762, n6496);
  and g12012 (n6497, n_5761, n_5762);
  and g12013 (n6498, n1666, n2334);
  and g12014 (n6499, n2115, n3110);
  and g12015 (n6500, n1919, n2617);
  not g12016 (n_5763, n6499);
  not g12017 (n_5764, n6500);
  and g12018 (n6501, n_5763, n_5764);
  not g12019 (n_5765, n6498);
  not g12020 (n_5766, n6501);
  and g12021 (n6502, n_5765, n_5766);
  not g12022 (n_5767, n6502);
  and g12023 (n6503, \a[30] , n_5767);
  and g12024 (n6504, \a[22] , n6503);
  and g12025 (n6505, \a[23] , \a[29] );
  and g12026 (n6506, \a[24] , \a[28] );
  not g12027 (n_5768, n6505);
  not g12028 (n_5769, n6506);
  and g12029 (n6507, n_5768, n_5769);
  and g12030 (n6508, n_5765, n_5767);
  not g12031 (n_5770, n6507);
  and g12032 (n6509, n_5770, n6508);
  not g12033 (n_5771, n6504);
  not g12034 (n_5772, n6509);
  and g12035 (n6510, n_5771, n_5772);
  not g12036 (n_5773, n6497);
  not g12037 (n_5774, n6510);
  and g12038 (n6511, n_5773, n_5774);
  not g12039 (n_5775, n6511);
  and g12040 (n6512, n_5773, n_5775);
  and g12041 (n6513, n_5774, n_5775);
  not g12042 (n_5776, n6512);
  not g12043 (n_5777, n6513);
  and g12044 (n6514, n_5776, n_5777);
  and g12045 (n6515, n5428, n6165);
  and g12046 (n6516, \a[9] , \a[43] );
  and g12047 (n6517, n4201, n6516);
  and g12048 (n6518, n745, n5083);
  not g12049 (n_5778, n6517);
  not g12050 (n_5779, n6518);
  and g12051 (n6519, n_5778, n_5779);
  not g12052 (n_5780, n6515);
  not g12053 (n_5781, n6519);
  and g12054 (n6520, n_5780, n_5781);
  not g12055 (n_5782, n6520);
  and g12056 (n6521, n4201, n_5782);
  and g12057 (n6522, n_5780, n_5782);
  and g12058 (n6523, \a[13] , \a[39] );
  not g12059 (n_5783, n6516);
  not g12060 (n_5784, n6523);
  and g12061 (n6524, n_5783, n_5784);
  not g12062 (n_5785, n6524);
  and g12063 (n6525, n6522, n_5785);
  not g12064 (n_5786, n6521);
  not g12065 (n_5787, n6525);
  and g12066 (n6526, n_5786, n_5787);
  not g12067 (n_5788, n6514);
  not g12068 (n_5789, n6526);
  and g12069 (n6527, n_5788, n_5789);
  not g12070 (n_5790, n6527);
  and g12071 (n6528, n_5788, n_5790);
  and g12072 (n6529, n_5789, n_5790);
  not g12073 (n_5791, n6528);
  not g12074 (n_5792, n6529);
  and g12075 (n6530, n_5791, n_5792);
  and g12076 (n6531, n6483, n6530);
  not g12077 (n_5793, n6483);
  not g12078 (n_5794, n6530);
  and g12079 (n6532, n_5793, n_5794);
  not g12080 (n_5795, n6531);
  not g12081 (n_5796, n6532);
  and g12082 (n6533, n_5795, n_5796);
  not g12083 (n_5797, n6436);
  and g12084 (n6534, n_5797, n6533);
  not g12085 (n_5798, n6533);
  and g12086 (n6535, n6436, n_5798);
  not g12087 (n_5799, n6534);
  not g12088 (n_5800, n6535);
  and g12089 (n6536, n_5799, n_5800);
  not g12090 (n_5801, n6435);
  and g12091 (n6537, n_5801, n6536);
  not g12092 (n_5802, n6536);
  and g12093 (n6538, n6435, n_5802);
  not g12094 (n_5803, n6537);
  not g12095 (n_5804, n6538);
  and g12096 (n6539, n_5803, n_5804);
  not g12097 (n_5805, n6539);
  and g12098 (n6540, n6434, n_5805);
  not g12099 (n_5806, n6434);
  and g12100 (n6541, n_5806, n6539);
  not g12101 (n_5807, n6540);
  not g12102 (n_5808, n6541);
  and g12103 (n6542, n_5807, n_5808);
  and g12104 (n6543, n_5529, n_5592);
  not g12105 (n_5809, n6543);
  and g12106 (n6544, n6542, n_5809);
  not g12107 (n_5810, n6542);
  and g12108 (n6545, n_5810, n6543);
  not g12109 (n_5811, n6544);
  not g12110 (n_5812, n6545);
  and g12111 (n6546, n_5811, n_5812);
  not g12112 (n_5813, n6433);
  and g12113 (n6547, n_5813, n6546);
  not g12114 (n_5814, n6546);
  and g12115 (n6548, n6433, n_5814);
  not g12116 (n_5815, n6547);
  not g12117 (n_5816, n6548);
  and g12118 (n6549, n_5815, n_5816);
  not g12119 (n_5817, n6549);
  and g12120 (n6550, n6319, n_5817);
  not g12121 (n_5818, n6319);
  and g12122 (n6551, n_5818, n6549);
  not g12123 (n_5819, n6550);
  not g12124 (n_5820, n6551);
  and g12125 (n6552, n_5819, n_5820);
  not g12126 (n_5821, n6552);
  and g12127 (n6553, n6318, n_5821);
  not g12128 (n_5822, n6318);
  and g12129 (n6554, n_5822, n_5819);
  and g12130 (n6555, n_5820, n6554);
  not g12131 (n_5823, n6553);
  not g12132 (n_5824, n6555);
  and g12133 (\asquared[53] , n_5823, n_5824);
  not g12134 (n_5825, n6554);
  and g12135 (n6557, n_5820, n_5825);
  and g12136 (n6558, n_5811, n_5815);
  and g12137 (n6559, n_5651, n_5713);
  and g12138 (n6560, n_5705, n_5709);
  and g12139 (n6561, \a[2] , \a[51] );
  and g12140 (n6562, \a[3] , \a[50] );
  not g12141 (n_5826, n6561);
  not g12142 (n_5827, n6562);
  and g12143 (n6563, n_5826, n_5827);
  and g12144 (n6564, \a[50] , \a[51] );
  and g12145 (n6565, n218, n6564);
  not g12146 (n_5828, n6563);
  not g12147 (n_5829, n6565);
  and g12148 (n6566, n_5828, n_5829);
  and g12149 (n6567, n6351, n6566);
  not g12150 (n_5830, n6567);
  and g12151 (n6568, n_5829, n_5830);
  and g12152 (n6569, n_5828, n6568);
  and g12153 (n6570, n6351, n_5830);
  not g12154 (n_5831, n6569);
  not g12155 (n_5832, n6570);
  and g12156 (n6571, n_5831, n_5832);
  and g12157 (n6572, \a[17] , \a[36] );
  and g12158 (n6573, \a[18] , \a[35] );
  not g12159 (n_5833, n6572);
  not g12160 (n_5834, n6573);
  and g12161 (n6574, n_5833, n_5834);
  and g12162 (n6575, n1052, n3828);
  not g12163 (n_5835, n6575);
  not g12166 (n_5836, n6574);
  not g12168 (n_5837, n6578);
  and g12169 (n6579, \a[49] , n_5837);
  and g12170 (n6580, \a[4] , n6579);
  and g12171 (n6581, n_5835, n_5837);
  and g12172 (n6582, n_5836, n6581);
  not g12173 (n_5838, n6580);
  not g12174 (n_5839, n6582);
  and g12175 (n6583, n_5838, n_5839);
  not g12176 (n_5840, n6571);
  not g12177 (n_5841, n6583);
  and g12178 (n6584, n_5840, n_5841);
  not g12179 (n_5842, n6584);
  and g12180 (n6585, n_5840, n_5842);
  and g12181 (n6586, n_5841, n_5842);
  not g12182 (n_5843, n6585);
  not g12183 (n_5844, n6586);
  and g12184 (n6587, n_5843, n_5844);
  and g12185 (n6588, n1494, n3143);
  and g12186 (n6589, n1492, n4090);
  and g12187 (n6590, n1490, n4150);
  not g12188 (n_5845, n6589);
  not g12189 (n_5846, n6590);
  and g12190 (n6591, n_5845, n_5846);
  not g12191 (n_5847, n6588);
  not g12192 (n_5848, n6591);
  and g12193 (n6592, n_5847, n_5848);
  not g12194 (n_5849, n6592);
  and g12195 (n6593, \a[34] , n_5849);
  and g12196 (n6594, \a[19] , n6593);
  and g12197 (n6595, n_5847, n_5849);
  and g12198 (n6596, \a[20] , \a[33] );
  and g12199 (n6597, \a[21] , \a[32] );
  not g12200 (n_5850, n6596);
  not g12201 (n_5851, n6597);
  and g12202 (n6598, n_5850, n_5851);
  not g12203 (n_5852, n6598);
  and g12204 (n6599, n6595, n_5852);
  not g12205 (n_5853, n6594);
  not g12206 (n_5854, n6599);
  and g12207 (n6600, n_5853, n_5854);
  not g12208 (n_5855, n6587);
  not g12209 (n_5856, n6600);
  and g12210 (n6601, n_5855, n_5856);
  not g12211 (n_5857, n6601);
  and g12212 (n6602, n_5855, n_5857);
  and g12213 (n6603, n_5856, n_5857);
  not g12214 (n_5858, n6602);
  not g12215 (n_5859, n6603);
  and g12216 (n6604, n_5858, n_5859);
  and g12217 (n6605, n_5614, n_5620);
  and g12218 (n6606, n6604, n6605);
  not g12219 (n_5860, n6604);
  not g12220 (n_5861, n6605);
  and g12221 (n6607, n_5860, n_5861);
  not g12222 (n_5862, n6606);
  not g12223 (n_5863, n6607);
  and g12224 (n6608, n_5862, n_5863);
  and g12225 (n6609, n335, n5666);
  and g12226 (n6610, \a[6] , \a[47] );
  and g12227 (n6611, n4204, n6610);
  not g12228 (n_5864, n6609);
  not g12229 (n_5865, n6611);
  and g12230 (n6612, n_5864, n_5865);
  and g12231 (n6613, \a[7] , \a[46] );
  and g12232 (n6614, n4204, n6613);
  not g12233 (n_5866, n6612);
  not g12234 (n_5867, n6614);
  and g12235 (n6615, n_5866, n_5867);
  not g12236 (n_5868, n6615);
  and g12237 (n6616, n_5867, n_5868);
  not g12238 (n_5869, n4204);
  not g12239 (n_5870, n6613);
  and g12240 (n6617, n_5869, n_5870);
  not g12241 (n_5871, n6617);
  and g12242 (n6618, n6616, n_5871);
  and g12243 (n6619, n6610, n_5868);
  not g12244 (n_5872, n6618);
  not g12245 (n_5873, n6619);
  and g12246 (n6620, n_5872, n_5873);
  and g12247 (n6621, \a[14] , \a[44] );
  and g12248 (n6622, n5428, n6621);
  and g12249 (n6623, n432, n5713);
  and g12250 (n6624, \a[8] , \a[45] );
  and g12251 (n6625, \a[14] , \a[39] );
  and g12252 (n6626, n6624, n6625);
  not g12253 (n_5874, n6623);
  not g12254 (n_5875, n6626);
  and g12255 (n6627, n_5874, n_5875);
  not g12256 (n_5876, n6622);
  not g12257 (n_5877, n6627);
  and g12258 (n6628, n_5876, n_5877);
  not g12259 (n_5878, n6628);
  and g12260 (n6629, n_5876, n_5878);
  and g12261 (n6630, \a[9] , \a[44] );
  not g12262 (n_5879, n6625);
  not g12263 (n_5880, n6630);
  and g12264 (n6631, n_5879, n_5880);
  not g12265 (n_5881, n6631);
  and g12266 (n6632, n6629, n_5881);
  and g12267 (n6633, n6624, n_5878);
  not g12268 (n_5882, n6632);
  not g12269 (n_5883, n6633);
  and g12270 (n6634, n_5882, n_5883);
  not g12271 (n_5884, n6620);
  not g12272 (n_5885, n6634);
  and g12273 (n6635, n_5884, n_5885);
  not g12274 (n_5886, n6635);
  and g12275 (n6636, n_5884, n_5886);
  and g12276 (n6637, n_5885, n_5886);
  not g12277 (n_5887, n6636);
  not g12278 (n_5888, n6637);
  and g12279 (n6638, n_5887, n_5888);
  and g12280 (n6639, \a[5] , \a[48] );
  and g12281 (n6640, \a[16] , \a[37] );
  not g12282 (n_5889, n6639);
  not g12283 (n_5890, n6640);
  and g12284 (n6641, n_5889, n_5890);
  and g12285 (n6642, \a[16] , \a[48] );
  and g12286 (n6643, n4242, n6642);
  not g12287 (n_5891, n6643);
  not g12290 (n_5893, n6641);
  not g12292 (n_5894, n6646);
  and g12293 (n6647, \a[53] , n_5894);
  and g12294 (n6648, \a[0] , n6647);
  and g12295 (n6649, n_5891, n_5894);
  and g12296 (n6650, n_5893, n6649);
  not g12297 (n_5895, n6648);
  not g12298 (n_5896, n6650);
  and g12299 (n6651, n_5895, n_5896);
  not g12300 (n_5897, n6638);
  not g12301 (n_5898, n6651);
  and g12302 (n6652, n_5897, n_5898);
  not g12303 (n_5899, n6652);
  and g12304 (n6653, n_5897, n_5899);
  and g12305 (n6654, n_5898, n_5899);
  not g12306 (n_5900, n6653);
  not g12307 (n_5901, n6654);
  and g12308 (n6655, n_5900, n_5901);
  not g12309 (n_5902, n6608);
  and g12310 (n6656, n_5902, n6655);
  not g12311 (n_5903, n6655);
  and g12312 (n6657, n6608, n_5903);
  not g12313 (n_5904, n6656);
  not g12314 (n_5905, n6657);
  and g12315 (n6658, n_5904, n_5905);
  and g12316 (n6659, \a[10] , \a[43] );
  and g12317 (n6660, \a[12] , \a[41] );
  not g12318 (n_5906, n6659);
  not g12319 (n_5907, n6660);
  and g12320 (n6661, n_5906, n_5907);
  and g12321 (n6662, n480, n4807);
  and g12322 (n6663, n5972, n6165);
  and g12323 (n6664, n748, n5413);
  not g12324 (n_5908, n6663);
  not g12325 (n_5909, n6664);
  and g12326 (n6665, n_5908, n_5909);
  not g12327 (n_5910, n6662);
  not g12328 (n_5911, n6665);
  and g12329 (n6666, n_5910, n_5911);
  not g12330 (n_5912, n6666);
  and g12331 (n6667, n_5910, n_5912);
  not g12332 (n_5913, n6661);
  and g12333 (n6668, n_5913, n6667);
  and g12334 (n6669, \a[40] , n_5912);
  and g12335 (n6670, \a[13] , n6669);
  not g12336 (n_5914, n6668);
  not g12337 (n_5915, n6670);
  and g12338 (n6671, n_5914, n_5915);
  and g12339 (n6672, n1666, n2617);
  and g12340 (n6673, n2115, n3452);
  and g12341 (n6674, n1919, n2865);
  not g12342 (n_5916, n6673);
  not g12343 (n_5917, n6674);
  and g12344 (n6675, n_5916, n_5917);
  not g12345 (n_5918, n6672);
  not g12346 (n_5919, n6675);
  and g12347 (n6676, n_5918, n_5919);
  not g12348 (n_5920, n6676);
  and g12349 (n6677, n2350, n_5920);
  and g12350 (n6678, \a[23] , \a[30] );
  and g12351 (n6679, \a[24] , \a[29] );
  not g12352 (n_5921, n6678);
  not g12353 (n_5922, n6679);
  and g12354 (n6680, n_5921, n_5922);
  and g12355 (n6681, n_5918, n_5920);
  not g12356 (n_5923, n6680);
  and g12357 (n6682, n_5923, n6681);
  not g12358 (n_5924, n6677);
  not g12359 (n_5925, n6682);
  and g12360 (n6683, n_5924, n_5925);
  not g12361 (n_5926, n6671);
  not g12362 (n_5927, n6683);
  and g12363 (n6684, n_5926, n_5927);
  not g12364 (n_5928, n6684);
  and g12365 (n6685, n_5926, n_5928);
  and g12366 (n6686, n_5927, n_5928);
  not g12367 (n_5929, n6685);
  not g12368 (n_5930, n6686);
  and g12369 (n6687, n_5929, n_5930);
  and g12370 (n6688, \a[25] , \a[28] );
  not g12371 (n_5931, n2227);
  not g12372 (n_5932, n6688);
  and g12373 (n6689, n_5931, n_5932);
  and g12374 (n6690, n2331, n2463);
  not g12375 (n_5933, n6690);
  not g12378 (n_5934, n6689);
  not g12380 (n_5935, n6693);
  and g12381 (n6694, \a[42] , n_5935);
  and g12382 (n6695, \a[11] , n6694);
  and g12383 (n6696, n_5933, n_5935);
  and g12384 (n6697, n_5934, n6696);
  not g12385 (n_5936, n6695);
  not g12386 (n_5937, n6697);
  and g12387 (n6698, n_5936, n_5937);
  not g12388 (n_5938, n6687);
  not g12389 (n_5939, n6698);
  and g12390 (n6699, n_5938, n_5939);
  not g12391 (n_5940, n6699);
  and g12392 (n6700, n_5938, n_5940);
  and g12393 (n6701, n_5939, n_5940);
  not g12394 (n_5941, n6700);
  not g12395 (n_5942, n6701);
  and g12396 (n6702, n_5941, n_5942);
  and g12397 (n6703, n_5638, n_5642);
  and g12398 (n6704, n6702, n6703);
  not g12399 (n_5943, n6702);
  not g12400 (n_5944, n6703);
  and g12401 (n6705, n_5943, n_5944);
  not g12402 (n_5945, n6704);
  not g12403 (n_5946, n6705);
  and g12404 (n6706, n_5945, n_5946);
  and g12405 (n6707, n_5699, n_5702);
  not g12406 (n_5947, n6707);
  and g12407 (n6708, n6706, n_5947);
  not g12408 (n_5948, n6706);
  and g12409 (n6709, n_5948, n6707);
  not g12410 (n_5949, n6708);
  not g12411 (n_5950, n6709);
  and g12412 (n6710, n_5949, n_5950);
  and g12413 (n6711, n6658, n6710);
  not g12414 (n_5951, n6658);
  not g12415 (n_5952, n6710);
  and g12416 (n6712, n_5951, n_5952);
  not g12417 (n_5953, n6711);
  not g12418 (n_5954, n6712);
  and g12419 (n6713, n_5953, n_5954);
  not g12420 (n_5955, n6560);
  and g12421 (n6714, n_5955, n6713);
  not g12422 (n_5956, n6713);
  and g12423 (n6715, n6560, n_5956);
  not g12424 (n_5957, n6714);
  not g12425 (n_5958, n6715);
  and g12426 (n6716, n_5957, n_5958);
  not g12427 (n_5959, n6559);
  and g12428 (n6717, n_5959, n6716);
  not g12429 (n_5960, n6716);
  and g12430 (n6718, n6559, n_5960);
  not g12431 (n_5961, n6717);
  not g12432 (n_5962, n6718);
  and g12433 (n6719, n_5961, n_5962);
  and g12434 (n6720, n6445, n6490);
  not g12435 (n_5963, n6445);
  not g12436 (n_5964, n6490);
  and g12437 (n6721, n_5963, n_5964);
  not g12438 (n_5965, n6720);
  not g12439 (n_5966, n6721);
  and g12440 (n6722, n_5965, n_5966);
  not g12441 (n_5967, n6722);
  and g12442 (n6723, n6477, n_5967);
  not g12443 (n_5968, n6477);
  and g12444 (n6724, n_5968, n6722);
  not g12445 (n_5969, n6723);
  not g12446 (n_5970, n6724);
  and g12447 (n6725, n_5969, n_5970);
  and g12448 (n6726, n_5738, n_5750);
  and g12449 (n6727, \a[52] , n1942);
  and g12450 (n6728, \a[1] , \a[52] );
  not g12451 (n_5971, \a[27] );
  not g12452 (n_5972, n6728);
  and g12453 (n6729, n_5971, n_5972);
  not g12454 (n_5973, n6727);
  not g12455 (n_5974, n6729);
  and g12456 (n6730, n_5973, n_5974);
  not g12457 (n_5975, n6730);
  and g12458 (n6731, n6459, n_5975);
  not g12459 (n_5976, n6459);
  and g12460 (n6732, n_5976, n6730);
  not g12461 (n_5977, n6731);
  not g12462 (n_5978, n6732);
  and g12463 (n6733, n_5977, n_5978);
  not g12464 (n_5979, n6522);
  and g12465 (n6734, n_5979, n6733);
  not g12466 (n_5980, n6733);
  and g12467 (n6735, n6522, n_5980);
  not g12468 (n_5981, n6734);
  not g12469 (n_5982, n6735);
  and g12470 (n6736, n_5981, n_5982);
  not g12471 (n_5983, n6726);
  and g12472 (n6737, n_5983, n6736);
  not g12473 (n_5984, n6737);
  and g12474 (n6738, n_5983, n_5984);
  and g12475 (n6739, n6736, n_5984);
  not g12476 (n_5985, n6738);
  not g12477 (n_5986, n6739);
  and g12478 (n6740, n_5985, n_5986);
  not g12479 (n_5987, n6740);
  and g12480 (n6741, n6725, n_5987);
  not g12481 (n_5988, n6741);
  and g12482 (n6742, n6725, n_5988);
  and g12483 (n6743, n_5987, n_5988);
  not g12484 (n_5989, n6742);
  not g12485 (n_5990, n6743);
  and g12486 (n6744, n_5989, n_5990);
  and g12487 (n6745, n6332, n6385);
  not g12488 (n_5991, n6332);
  not g12489 (n_5992, n6385);
  and g12490 (n6746, n_5991, n_5992);
  not g12491 (n_5993, n6745);
  not g12492 (n_5994, n6746);
  and g12493 (n6747, n_5993, n_5994);
  not g12494 (n_5995, n6747);
  and g12495 (n6748, n6508, n_5995);
  not g12496 (n_5996, n6508);
  and g12497 (n6749, n_5996, n6747);
  not g12498 (n_5997, n6748);
  not g12499 (n_5998, n6749);
  and g12500 (n6750, n_5997, n_5998);
  and g12501 (n6751, n_5775, n_5790);
  and g12502 (n6752, n_5655, n_5668);
  and g12503 (n6753, n6751, n6752);
  not g12504 (n_5999, n6751);
  not g12505 (n_6000, n6752);
  and g12506 (n6754, n_5999, n_6000);
  not g12507 (n_6001, n6753);
  not g12508 (n_6002, n6754);
  and g12509 (n6755, n_6001, n_6002);
  and g12510 (n6756, n6750, n6755);
  not g12511 (n_6003, n6750);
  not g12512 (n_6004, n6755);
  and g12513 (n6757, n_6003, n_6004);
  not g12514 (n_6005, n6756);
  not g12515 (n_6006, n6757);
  and g12516 (n6758, n_6005, n_6006);
  not g12517 (n_6007, n6744);
  and g12518 (n6759, n_6007, n6758);
  not g12519 (n_6008, n6759);
  and g12520 (n6760, n6758, n_6008);
  and g12521 (n6761, n_6007, n_6008);
  not g12522 (n_6009, n6760);
  not g12523 (n_6010, n6761);
  and g12524 (n6762, n_6009, n_6010);
  and g12525 (n6763, n_5624, n_5646);
  and g12526 (n6764, n6762, n6763);
  not g12527 (n_6011, n6762);
  not g12528 (n_6012, n6763);
  and g12529 (n6765, n_6011, n_6012);
  not g12530 (n_6013, n6764);
  not g12531 (n_6014, n6765);
  and g12532 (n6766, n_6013, n_6014);
  and g12533 (n6767, n_5796, n_5799);
  and g12534 (n6768, n_5683, n_5687);
  and g12535 (n6769, n_5630, n_5634);
  and g12536 (n6770, n6768, n6769);
  not g12537 (n_6015, n6768);
  not g12538 (n_6016, n6769);
  and g12539 (n6771, n_6015, n_6016);
  not g12540 (n_6017, n6770);
  not g12541 (n_6018, n6771);
  and g12542 (n6772, n_6017, n_6018);
  and g12543 (n6773, n_5691, n_5695);
  not g12544 (n_6019, n6772);
  and g12545 (n6774, n_6019, n6773);
  not g12546 (n_6020, n6773);
  and g12547 (n6775, n6772, n_6020);
  not g12548 (n_6021, n6774);
  not g12549 (n_6022, n6775);
  and g12550 (n6776, n_6021, n_6022);
  and g12551 (n6777, n_5674, n_5678);
  not g12552 (n_6023, n6776);
  and g12553 (n6778, n_6023, n6777);
  not g12554 (n_6024, n6777);
  and g12555 (n6779, n6776, n_6024);
  not g12556 (n_6025, n6778);
  not g12557 (n_6026, n6779);
  and g12558 (n6780, n_6025, n_6026);
  not g12559 (n_6027, n6767);
  and g12560 (n6781, n_6027, n6780);
  not g12561 (n_6028, n6780);
  and g12562 (n6782, n6767, n_6028);
  not g12563 (n_6029, n6781);
  not g12564 (n_6030, n6782);
  and g12565 (n6783, n_6029, n_6030);
  and g12566 (n6784, n_5803, n_5808);
  not g12567 (n_6031, n6783);
  and g12568 (n6785, n_6031, n6784);
  not g12569 (n_6032, n6784);
  and g12570 (n6786, n6783, n_6032);
  not g12571 (n_6033, n6785);
  not g12572 (n_6034, n6786);
  and g12573 (n6787, n_6033, n_6034);
  and g12574 (n6788, n6766, n6787);
  not g12575 (n_6035, n6766);
  not g12576 (n_6036, n6787);
  and g12577 (n6789, n_6035, n_6036);
  not g12578 (n_6037, n6788);
  not g12579 (n_6038, n6789);
  and g12580 (n6790, n_6037, n_6038);
  and g12581 (n6791, n6719, n6790);
  not g12582 (n_6039, n6719);
  not g12583 (n_6040, n6790);
  and g12584 (n6792, n_6039, n_6040);
  not g12585 (n_6041, n6791);
  not g12586 (n_6042, n6792);
  and g12587 (n6793, n_6041, n_6042);
  not g12588 (n_6043, n6558);
  and g12589 (n6794, n_6043, n6793);
  not g12590 (n_6044, n6793);
  and g12591 (n6795, n6558, n_6044);
  not g12592 (n_6045, n6794);
  not g12593 (n_6046, n6795);
  and g12594 (n6796, n_6045, n_6046);
  not g12595 (n_6047, n6557);
  not g12596 (n_6048, n6796);
  and g12597 (n6797, n_6047, n_6048);
  and g12598 (n6798, n6557, n6796);
  or g12599 (\asquared[54] , n6797, n6798);
  and g12600 (n6800, n_5961, n_6041);
  and g12601 (n6801, n_6008, n_6014);
  and g12602 (n6802, n_6026, n_6029);
  and g12603 (n6803, n6801, n6802);
  not g12604 (n_6049, n6801);
  not g12605 (n_6050, n6802);
  and g12606 (n6804, n_6049, n_6050);
  not g12607 (n_6051, n6803);
  not g12608 (n_6052, n6804);
  and g12609 (n6805, n_6051, n_6052);
  and g12610 (n6806, n_5984, n_5988);
  and g12611 (n6807, n_6002, n_6005);
  and g12612 (n6808, \a[0] , \a[54] );
  and g12613 (n6809, n6727, n6808);
  not g12614 (n_6054, n6809);
  and g12615 (n6810, n6727, n_6054);
  and g12616 (n6811, n_5973, n6808);
  not g12617 (n_6055, n6810);
  not g12618 (n_6056, n6811);
  and g12619 (n6812, n_6055, n_6056);
  and g12620 (n6813, \a[1] , \a[53] );
  and g12621 (n6814, n2800, n6813);
  not g12622 (n_6057, n6814);
  and g12623 (n6815, n6813, n_6057);
  and g12624 (n6816, n2800, n_6057);
  not g12625 (n_6058, n6815);
  not g12626 (n_6059, n6816);
  and g12627 (n6817, n_6058, n_6059);
  not g12628 (n_6060, n6812);
  not g12629 (n_6061, n6817);
  and g12630 (n6818, n_6060, n_6061);
  not g12631 (n_6062, n6818);
  and g12632 (n6819, n_6060, n_6062);
  and g12633 (n6820, n_6061, n_6062);
  not g12634 (n_6063, n6819);
  not g12635 (n_6064, n6820);
  and g12636 (n6821, n_6063, n_6064);
  and g12637 (n6822, n1574, n3143);
  and g12638 (n6823, \a[32] , \a[35] );
  and g12639 (n6824, n4036, n6823);
  and g12640 (n6825, n1492, n2972);
  not g12641 (n_6065, n6824);
  not g12642 (n_6066, n6825);
  and g12643 (n6826, n_6065, n_6066);
  not g12644 (n_6067, n6822);
  not g12645 (n_6068, n6826);
  and g12646 (n6827, n_6067, n_6068);
  not g12647 (n_6069, n6827);
  and g12648 (n6828, n_6067, n_6069);
  and g12649 (n6829, \a[21] , \a[33] );
  and g12650 (n6830, \a[22] , \a[32] );
  not g12651 (n_6070, n6829);
  not g12652 (n_6071, n6830);
  and g12653 (n6831, n_6070, n_6071);
  not g12654 (n_6072, n6831);
  and g12655 (n6832, n6828, n_6072);
  and g12656 (n6833, \a[35] , n_6069);
  and g12657 (n6834, \a[19] , n6833);
  not g12658 (n_6073, n6832);
  not g12659 (n_6074, n6834);
  and g12660 (n6835, n_6073, n_6074);
  and g12661 (n6836, n1904, n2617);
  and g12662 (n6837, n1547, n3452);
  and g12663 (n6838, n1666, n2865);
  not g12664 (n_6075, n6837);
  not g12665 (n_6076, n6838);
  and g12666 (n6839, n_6075, n_6076);
  not g12667 (n_6077, n6836);
  not g12668 (n_6078, n6839);
  and g12669 (n6840, n_6077, n_6078);
  not g12670 (n_6079, n6840);
  and g12671 (n6841, \a[31] , n_6079);
  and g12672 (n6842, \a[23] , n6841);
  and g12673 (n6843, n_6077, n_6079);
  and g12674 (n6844, \a[25] , \a[29] );
  not g12675 (n_6080, n2619);
  not g12676 (n_6081, n6844);
  and g12677 (n6845, n_6080, n_6081);
  not g12678 (n_6082, n6845);
  and g12679 (n6846, n6843, n_6082);
  not g12680 (n_6083, n6842);
  not g12681 (n_6084, n6846);
  and g12682 (n6847, n_6083, n_6084);
  not g12683 (n_6085, n6835);
  not g12684 (n_6086, n6847);
  and g12685 (n6848, n_6085, n_6086);
  not g12686 (n_6087, n6848);
  and g12687 (n6849, n_6085, n_6087);
  and g12688 (n6850, n_6086, n_6087);
  not g12689 (n_6088, n6849);
  not g12690 (n_6089, n6850);
  and g12691 (n6851, n_6088, n_6089);
  not g12692 (n_6090, n6821);
  and g12693 (n6852, n_6090, n6851);
  not g12694 (n_6091, n6851);
  and g12695 (n6853, n6821, n_6091);
  not g12696 (n_6092, n6852);
  not g12697 (n_6093, n6853);
  and g12698 (n6854, n_6092, n_6093);
  not g12699 (n_6094, n6807);
  not g12700 (n_6095, n6854);
  and g12701 (n6855, n_6094, n_6095);
  not g12702 (n_6096, n6855);
  and g12703 (n6856, n_6094, n_6096);
  and g12704 (n6857, n_6095, n_6096);
  not g12705 (n_6097, n6856);
  not g12706 (n_6098, n6857);
  and g12707 (n6858, n_6097, n_6098);
  not g12708 (n_6099, n6806);
  not g12709 (n_6100, n6858);
  and g12710 (n6859, n_6099, n_6100);
  not g12711 (n_6101, n6859);
  and g12712 (n6860, n_6099, n_6101);
  and g12713 (n6861, n_6100, n_6101);
  not g12714 (n_6102, n6860);
  not g12715 (n_6103, n6861);
  and g12716 (n6862, n_6102, n_6103);
  not g12717 (n_6104, n6862);
  and g12718 (n6863, n6805, n_6104);
  not g12719 (n_6105, n6863);
  and g12720 (n6864, n6805, n_6105);
  and g12721 (n6865, n_6104, n_6105);
  not g12722 (n_6106, n6864);
  not g12723 (n_6107, n6865);
  and g12724 (n6866, n_6106, n_6107);
  and g12725 (n6867, n_6034, n_6037);
  not g12726 (n_6108, n6866);
  not g12727 (n_6109, n6867);
  and g12728 (n6868, n_6108, n_6109);
  not g12729 (n_6110, n6868);
  and g12730 (n6869, n_6108, n_6110);
  and g12731 (n6870, n_6109, n_6110);
  not g12732 (n_6111, n6869);
  not g12733 (n_6112, n6870);
  and g12734 (n6871, n_6111, n_6112);
  and g12735 (n6872, n_5953, n_5957);
  and g12736 (n6873, n_5966, n_5970);
  and g12737 (n6874, n_5994, n_5998);
  and g12738 (n6875, n6873, n6874);
  not g12739 (n_6113, n6873);
  not g12740 (n_6114, n6874);
  and g12741 (n6876, n_6113, n_6114);
  not g12742 (n_6115, n6875);
  not g12743 (n_6116, n6876);
  and g12744 (n6877, n_6115, n_6116);
  and g12745 (n6878, n_5978, n_5981);
  not g12746 (n_6117, n6877);
  and g12747 (n6879, n_6117, n6878);
  not g12748 (n_6118, n6878);
  and g12749 (n6880, n6877, n_6118);
  not g12750 (n_6119, n6879);
  not g12751 (n_6120, n6880);
  and g12752 (n6881, n_6119, n_6120);
  and g12753 (n6882, n_5863, n_5905);
  not g12754 (n_6121, n6882);
  and g12755 (n6883, n6881, n_6121);
  not g12756 (n_6122, n6881);
  and g12757 (n6884, n_6122, n6882);
  not g12758 (n_6123, n6883);
  not g12759 (n_6124, n6884);
  and g12760 (n6885, n_6123, n_6124);
  and g12761 (n6886, n6616, n6649);
  not g12762 (n_6125, n6616);
  not g12763 (n_6126, n6649);
  and g12764 (n6887, n_6125, n_6126);
  not g12765 (n_6127, n6886);
  not g12766 (n_6128, n6887);
  and g12767 (n6888, n_6127, n_6128);
  not g12768 (n_6129, n6888);
  and g12769 (n6889, n6696, n_6129);
  not g12770 (n_6130, n6696);
  and g12771 (n6890, n_6130, n6888);
  not g12772 (n_6131, n6889);
  not g12773 (n_6132, n6890);
  and g12774 (n6891, n_6131, n_6132);
  and g12775 (n6892, n6581, n6595);
  not g12776 (n_6133, n6581);
  not g12777 (n_6134, n6595);
  and g12778 (n6893, n_6133, n_6134);
  not g12779 (n_6135, n6892);
  not g12780 (n_6136, n6893);
  and g12781 (n6894, n_6135, n_6136);
  not g12782 (n_6137, n6894);
  and g12783 (n6895, n6681, n_6137);
  not g12784 (n_6138, n6681);
  and g12785 (n6896, n_6138, n6894);
  not g12786 (n_6139, n6895);
  not g12787 (n_6140, n6896);
  and g12788 (n6897, n_6139, n_6140);
  and g12789 (n6898, n_5886, n_5899);
  not g12790 (n_6141, n6897);
  and g12791 (n6899, n_6141, n6898);
  not g12792 (n_6142, n6898);
  and g12793 (n6900, n6897, n_6142);
  not g12794 (n_6143, n6899);
  not g12795 (n_6144, n6900);
  and g12796 (n6901, n_6143, n_6144);
  and g12797 (n6902, n6891, n6901);
  not g12798 (n_6145, n6891);
  not g12799 (n_6146, n6901);
  and g12800 (n6903, n_6145, n_6146);
  not g12801 (n_6147, n6902);
  not g12802 (n_6148, n6903);
  and g12803 (n6904, n_6147, n_6148);
  and g12804 (n6905, n6885, n6904);
  not g12805 (n_6149, n6885);
  not g12806 (n_6150, n6904);
  and g12807 (n6906, n_6149, n_6150);
  not g12808 (n_6151, n6905);
  not g12809 (n_6152, n6906);
  and g12810 (n6907, n_6151, n_6152);
  not g12811 (n_6153, n6907);
  and g12812 (n6908, n6872, n_6153);
  not g12813 (n_6154, n6872);
  and g12814 (n6909, n_6154, n6907);
  not g12815 (n_6155, n6908);
  not g12816 (n_6156, n6909);
  and g12817 (n6910, n_6155, n_6156);
  and g12818 (n6911, \a[5] , \a[49] );
  and g12819 (n6912, \a[18] , \a[36] );
  not g12820 (n_6157, n6911);
  not g12821 (n_6158, n6912);
  and g12822 (n6913, n_6157, n_6158);
  and g12823 (n6914, \a[20] , \a[49] );
  and g12824 (n6915, n3664, n6914);
  and g12825 (n6916, n1331, n4595);
  not g12826 (n_6159, n6915);
  not g12827 (n_6160, n6916);
  and g12828 (n6917, n_6159, n_6160);
  and g12829 (n6918, n6911, n6912);
  not g12830 (n_6161, n6917);
  not g12831 (n_6162, n6918);
  and g12832 (n6919, n_6161, n_6162);
  not g12833 (n_6163, n6919);
  and g12834 (n6920, n_6162, n_6163);
  not g12835 (n_6164, n6913);
  and g12836 (n6921, n_6164, n6920);
  and g12837 (n6922, \a[34] , n_6163);
  and g12838 (n6923, \a[20] , n6922);
  not g12839 (n_6165, n6921);
  not g12840 (n_6166, n6923);
  and g12841 (n6924, n_6165, n_6166);
  and g12842 (n6925, n602, n5018);
  and g12843 (n6926, n818, n4807);
  and g12844 (n6927, n748, n5344);
  not g12845 (n_6167, n6926);
  not g12846 (n_6168, n6927);
  and g12847 (n6928, n_6167, n_6168);
  not g12848 (n_6169, n6925);
  not g12849 (n_6170, n6928);
  and g12850 (n6929, n_6169, n_6170);
  not g12851 (n_6171, n6929);
  and g12852 (n6930, \a[41] , n_6171);
  and g12853 (n6931, \a[13] , n6930);
  and g12854 (n6932, n_6169, n_6171);
  and g12855 (n6933, \a[11] , \a[43] );
  and g12856 (n6934, \a[12] , \a[42] );
  not g12857 (n_6172, n6933);
  not g12858 (n_6173, n6934);
  and g12859 (n6935, n_6172, n_6173);
  not g12860 (n_6174, n6935);
  and g12861 (n6936, n6932, n_6174);
  not g12862 (n_6175, n6931);
  not g12863 (n_6176, n6936);
  and g12864 (n6937, n_6175, n_6176);
  not g12865 (n_6177, n6924);
  not g12866 (n_6178, n6937);
  and g12867 (n6938, n_6177, n_6178);
  not g12868 (n_6179, n6938);
  and g12869 (n6939, n_6177, n_6179);
  and g12870 (n6940, n_6178, n_6179);
  not g12871 (n_6180, n6939);
  not g12872 (n_6181, n6940);
  and g12873 (n6941, n_6180, n_6181);
  and g12874 (n6942, \a[38] , \a[48] );
  and g12875 (n6943, n721, n6942);
  and g12876 (n6944, \a[17] , \a[48] );
  and g12877 (n6945, n4488, n6944);
  and g12878 (n6946, n1048, n4565);
  not g12879 (n_6182, n6945);
  not g12880 (n_6183, n6946);
  and g12881 (n6947, n_6182, n_6183);
  not g12882 (n_6184, n6943);
  not g12883 (n_6185, n6947);
  and g12884 (n6948, n_6184, n_6185);
  not g12885 (n_6186, n6948);
  and g12886 (n6949, \a[37] , n_6186);
  and g12887 (n6950, \a[17] , n6949);
  and g12888 (n6951, \a[6] , \a[48] );
  and g12889 (n6952, \a[16] , \a[38] );
  not g12890 (n_6187, n6951);
  not g12891 (n_6188, n6952);
  and g12892 (n6953, n_6187, n_6188);
  and g12893 (n6954, n_6184, n_6186);
  not g12894 (n_6189, n6953);
  and g12895 (n6955, n_6189, n6954);
  not g12896 (n_6190, n6950);
  not g12897 (n_6191, n6955);
  and g12898 (n6956, n_6190, n_6191);
  not g12899 (n_6192, n6941);
  not g12900 (n_6193, n6956);
  and g12901 (n6957, n_6192, n_6193);
  not g12902 (n_6194, n6957);
  and g12903 (n6958, n_6192, n_6194);
  and g12904 (n6959, n_6193, n_6194);
  not g12905 (n_6195, n6958);
  not g12906 (n_6196, n6959);
  and g12907 (n6960, n_6195, n_6196);
  and g12908 (n6961, n_6018, n_6022);
  and g12909 (n6962, n6960, n6961);
  not g12910 (n_6197, n6960);
  not g12911 (n_6198, n6961);
  and g12912 (n6963, n_6197, n_6198);
  not g12913 (n_6199, n6962);
  not g12914 (n_6200, n6963);
  and g12915 (n6964, n_6199, n_6200);
  and g12916 (n6965, n209, n6564);
  and g12917 (n6966, \a[50] , \a[52] );
  and g12918 (n6967, n252, n6966);
  and g12919 (n6968, \a[51] , \a[52] );
  and g12920 (n6969, n218, n6968);
  not g12921 (n_6201, n6967);
  not g12922 (n_6202, n6969);
  and g12923 (n6970, n_6201, n_6202);
  not g12924 (n_6203, n6965);
  not g12925 (n_6204, n6970);
  and g12926 (n6971, n_6203, n_6204);
  not g12927 (n_6205, n6971);
  and g12928 (n6972, n_6203, n_6205);
  and g12929 (n6973, \a[3] , \a[51] );
  and g12930 (n6974, \a[4] , \a[50] );
  not g12931 (n_6206, n6973);
  not g12932 (n_6207, n6974);
  and g12933 (n6975, n_6206, n_6207);
  not g12934 (n_6208, n6975);
  and g12935 (n6976, n6972, n_6208);
  and g12936 (n6977, \a[52] , n_6205);
  and g12937 (n6978, \a[2] , n6977);
  not g12938 (n_6209, n6976);
  not g12939 (n_6210, n6978);
  and g12940 (n6979, n_6209, n_6210);
  and g12941 (n6980, \a[7] , \a[47] );
  and g12942 (n6981, \a[15] , \a[39] );
  and g12943 (n6982, n6980, n6981);
  and g12944 (n6983, n380, n5666);
  not g12945 (n_6211, n6982);
  not g12946 (n_6212, n6983);
  and g12947 (n6984, n_6211, n_6212);
  and g12948 (n6985, \a[8] , \a[46] );
  and g12949 (n6986, n6981, n6985);
  not g12950 (n_6213, n6984);
  not g12951 (n_6214, n6986);
  and g12952 (n6987, n_6213, n_6214);
  not g12953 (n_6215, n6987);
  and g12954 (n6988, n6980, n_6215);
  and g12955 (n6989, n_6214, n_6215);
  not g12956 (n_6216, n6981);
  not g12957 (n_6217, n6985);
  and g12958 (n6990, n_6216, n_6217);
  not g12959 (n_6218, n6990);
  and g12960 (n6991, n6989, n_6218);
  not g12961 (n_6219, n6988);
  not g12962 (n_6220, n6991);
  and g12963 (n6992, n_6219, n_6220);
  not g12964 (n_6221, n6979);
  not g12965 (n_6222, n6992);
  and g12966 (n6993, n_6221, n_6222);
  not g12967 (n_6223, n6993);
  and g12968 (n6994, n_6221, n_6223);
  and g12969 (n6995, n_6222, n_6223);
  not g12970 (n_6224, n6994);
  not g12971 (n_6225, n6995);
  and g12972 (n6996, n_6224, n_6225);
  and g12973 (n6997, \a[9] , \a[45] );
  and g12974 (n6998, n5972, n6621);
  and g12975 (n6999, n484, n5713);
  and g12976 (n7000, n4855, n6997);
  not g12977 (n_6226, n6999);
  not g12978 (n_6227, n7000);
  and g12979 (n7001, n_6226, n_6227);
  not g12980 (n_6228, n6998);
  not g12981 (n_6229, n7001);
  and g12982 (n7002, n_6228, n_6229);
  not g12983 (n_6230, n7002);
  and g12984 (n7003, n6997, n_6230);
  and g12985 (n7004, n_6228, n_6230);
  and g12986 (n7005, \a[10] , \a[44] );
  not g12987 (n_6231, n4855);
  not g12988 (n_6232, n7005);
  and g12989 (n7006, n_6231, n_6232);
  not g12990 (n_6233, n7006);
  and g12991 (n7007, n7004, n_6233);
  not g12992 (n_6234, n7003);
  not g12993 (n_6235, n7007);
  and g12994 (n7008, n_6234, n_6235);
  not g12995 (n_6236, n6996);
  not g12996 (n_6237, n7008);
  and g12997 (n7009, n_6236, n_6237);
  not g12998 (n_6238, n7009);
  and g12999 (n7010, n_6236, n_6238);
  and g13000 (n7011, n_6237, n_6238);
  not g13001 (n_6239, n7010);
  not g13002 (n_6240, n7011);
  and g13003 (n7012, n_6239, n_6240);
  not g13004 (n_6241, n6964);
  and g13005 (n7013, n_6241, n7012);
  not g13006 (n_6242, n7012);
  and g13007 (n7014, n6964, n_6242);
  not g13008 (n_6243, n7013);
  not g13009 (n_6244, n7014);
  and g13010 (n7015, n_6243, n_6244);
  and g13011 (n7016, n_5946, n_5949);
  and g13012 (n7017, n6568, n6629);
  not g13013 (n_6245, n6568);
  not g13014 (n_6246, n6629);
  and g13015 (n7018, n_6245, n_6246);
  not g13016 (n_6247, n7017);
  not g13017 (n_6248, n7018);
  and g13018 (n7019, n_6247, n_6248);
  not g13019 (n_6249, n7019);
  and g13020 (n7020, n6667, n_6249);
  not g13021 (n_6250, n6667);
  and g13022 (n7021, n_6250, n7019);
  not g13023 (n_6251, n7020);
  not g13024 (n_6252, n7021);
  and g13025 (n7022, n_6251, n_6252);
  and g13026 (n7023, n_5928, n_5940);
  and g13027 (n7024, n_5842, n_5857);
  and g13028 (n7025, n7023, n7024);
  not g13029 (n_6253, n7023);
  not g13030 (n_6254, n7024);
  and g13031 (n7026, n_6253, n_6254);
  not g13032 (n_6255, n7025);
  not g13033 (n_6256, n7026);
  and g13034 (n7027, n_6255, n_6256);
  and g13035 (n7028, n7022, n7027);
  not g13036 (n_6257, n7022);
  not g13037 (n_6258, n7027);
  and g13038 (n7029, n_6257, n_6258);
  not g13039 (n_6259, n7028);
  not g13040 (n_6260, n7029);
  and g13041 (n7030, n_6259, n_6260);
  not g13042 (n_6261, n7016);
  and g13043 (n7031, n_6261, n7030);
  not g13044 (n_6262, n7031);
  and g13045 (n7032, n_6261, n_6262);
  and g13046 (n7033, n7030, n_6262);
  not g13047 (n_6263, n7032);
  not g13048 (n_6264, n7033);
  and g13049 (n7034, n_6263, n_6264);
  not g13050 (n_6265, n7034);
  and g13051 (n7035, n7015, n_6265);
  not g13052 (n_6266, n7035);
  and g13053 (n7036, n7015, n_6266);
  and g13054 (n7037, n_6265, n_6266);
  not g13055 (n_6267, n7036);
  not g13056 (n_6268, n7037);
  and g13057 (n7038, n_6267, n_6268);
  not g13058 (n_6269, n7038);
  and g13059 (n7039, n6910, n_6269);
  not g13060 (n_6270, n7039);
  and g13061 (n7040, n6910, n_6270);
  and g13062 (n7041, n_6269, n_6270);
  not g13063 (n_6271, n7040);
  not g13064 (n_6272, n7041);
  and g13065 (n7042, n_6271, n_6272);
  not g13066 (n_6273, n6871);
  and g13067 (n7043, n_6273, n7042);
  not g13068 (n_6274, n7042);
  and g13069 (n7044, n6871, n_6274);
  not g13070 (n_6275, n7043);
  not g13071 (n_6276, n7044);
  and g13072 (n7045, n_6275, n_6276);
  not g13073 (n_6277, n6800);
  not g13074 (n_6278, n7045);
  and g13075 (n7046, n_6277, n_6278);
  and g13076 (n7047, n6800, n7045);
  not g13077 (n_6279, n7046);
  not g13078 (n_6280, n7047);
  and g13079 (n7048, n_6279, n_6280);
  and g13080 (n7049, n_6047, n_6046);
  not g13081 (n_6281, n7049);
  and g13082 (n7050, n_6045, n_6281);
  not g13083 (n_6282, n7048);
  and g13084 (n7051, n_6282, n7050);
  not g13085 (n_6283, n7050);
  and g13086 (n7052, n7048, n_6283);
  not g13087 (n_6284, n7051);
  not g13088 (n_6285, n7052);
  and g13089 (\asquared[55] , n_6284, n_6285);
  and g13090 (n7054, n_6273, n_6274);
  not g13091 (n_6286, n7054);
  and g13092 (n7055, n_6110, n_6286);
  and g13093 (n7056, n_6156, n_6270);
  and g13094 (n7057, n_6262, n_6266);
  and g13095 (n7058, n_6123, n_6151);
  and g13096 (n7059, n_6144, n_6147);
  and g13097 (n7060, \a[6] , \a[49] );
  and g13098 (n7061, \a[17] , \a[38] );
  not g13099 (n_6287, n7060);
  not g13100 (n_6288, n7061);
  and g13101 (n7062, n_6287, n_6288);
  and g13102 (n7063, \a[17] , \a[49] );
  and g13103 (n7064, n4560, n7063);
  not g13104 (n_6289, n7064);
  not g13107 (n_6290, n7062);
  not g13109 (n_6291, n7067);
  and g13110 (n7068, n_6289, n_6291);
  and g13111 (n7069, n_6290, n7068);
  and g13112 (n7070, \a[52] , n_6291);
  and g13113 (n7071, \a[3] , n7070);
  not g13114 (n_6292, n7069);
  not g13115 (n_6293, n7071);
  and g13116 (n7072, n_6292, n_6293);
  and g13117 (n7073, \a[40] , \a[46] );
  and g13118 (n7074, n1517, n7073);
  and g13119 (n7075, n895, n5413);
  not g13120 (n_6294, n7074);
  not g13121 (n_6295, n7075);
  and g13122 (n7076, n_6294, n_6295);
  and g13123 (n7077, \a[9] , \a[46] );
  and g13124 (n7078, \a[14] , \a[41] );
  and g13125 (n7079, n7077, n7078);
  not g13126 (n_6296, n7076);
  not g13127 (n_6297, n7079);
  and g13128 (n7080, n_6296, n_6297);
  not g13129 (n_6298, n7080);
  and g13130 (n7081, \a[40] , n_6298);
  and g13131 (n7082, \a[15] , n7081);
  not g13132 (n_6299, n7077);
  not g13133 (n_6300, n7078);
  and g13134 (n7083, n_6299, n_6300);
  and g13135 (n7084, n_6297, n_6298);
  not g13136 (n_6301, n7083);
  and g13137 (n7085, n_6301, n7084);
  not g13138 (n_6302, n7082);
  not g13139 (n_6303, n7085);
  and g13140 (n7086, n_6302, n_6303);
  not g13141 (n_6304, n7072);
  not g13142 (n_6305, n7086);
  and g13143 (n7087, n_6304, n_6305);
  not g13144 (n_6306, n7087);
  and g13145 (n7088, n_6304, n_6306);
  and g13146 (n7089, n_6305, n_6306);
  not g13147 (n_6307, n7088);
  not g13148 (n_6308, n7089);
  and g13149 (n7090, n_6307, n_6308);
  and g13150 (n7091, n_6136, n_6140);
  and g13151 (n7092, n7090, n7091);
  not g13152 (n_6309, n7090);
  not g13153 (n_6310, n7091);
  and g13154 (n7093, n_6309, n_6310);
  not g13155 (n_6311, n7092);
  not g13156 (n_6312, n7093);
  and g13157 (n7094, n_6311, n_6312);
  and g13158 (n7095, n_6256, n_6259);
  not g13159 (n_6313, n7095);
  and g13160 (n7096, n7094, n_6313);
  not g13161 (n_6314, n7094);
  and g13162 (n7097, n_6314, n7095);
  not g13163 (n_6315, n7096);
  not g13164 (n_6316, n7097);
  and g13165 (n7098, n_6315, n_6316);
  not g13166 (n_6317, n7059);
  and g13167 (n7099, n_6317, n7098);
  not g13168 (n_6318, n7098);
  and g13169 (n7100, n7059, n_6318);
  not g13170 (n_6319, n7099);
  not g13171 (n_6320, n7100);
  and g13172 (n7101, n_6319, n_6320);
  not g13173 (n_6321, n7058);
  and g13174 (n7102, n_6321, n7101);
  not g13175 (n_6322, n7102);
  and g13176 (n7103, n_6321, n_6322);
  and g13177 (n7104, n7101, n_6322);
  not g13178 (n_6323, n7103);
  not g13179 (n_6324, n7104);
  and g13180 (n7105, n_6323, n_6324);
  not g13181 (n_6325, n7057);
  not g13182 (n_6326, n7105);
  and g13183 (n7106, n_6325, n_6326);
  not g13184 (n_6327, n7106);
  and g13185 (n7107, n_6325, n_6327);
  and g13186 (n7108, n_6326, n_6327);
  not g13187 (n_6328, n7107);
  not g13188 (n_6329, n7108);
  and g13189 (n7109, n_6328, n_6329);
  not g13190 (n_6330, n7056);
  not g13191 (n_6331, n7109);
  and g13192 (n7110, n_6330, n_6331);
  not g13193 (n_6332, n7110);
  and g13194 (n7111, n_6330, n_6332);
  and g13195 (n7112, n_6331, n_6332);
  not g13196 (n_6333, n7111);
  not g13197 (n_6334, n7112);
  and g13198 (n7113, n_6333, n_6334);
  and g13199 (n7114, n_6128, n_6132);
  and g13200 (n7115, n_6248, n_6252);
  and g13201 (n7116, n7114, n7115);
  not g13202 (n_6335, n7114);
  not g13203 (n_6336, n7115);
  and g13204 (n7117, n_6335, n_6336);
  not g13205 (n_6337, n7116);
  not g13206 (n_6338, n7117);
  and g13207 (n7118, n_6337, n_6338);
  and g13208 (n7119, \a[28] , \a[54] );
  and g13209 (n7120, \a[1] , n7119);
  and g13210 (n7121, \a[1] , \a[54] );
  not g13211 (n_6339, \a[28] );
  not g13212 (n_6340, n7121);
  and g13213 (n7122, n_6339, n_6340);
  not g13214 (n_6341, n7120);
  not g13215 (n_6342, n7122);
  and g13216 (n7123, n_6341, n_6342);
  and g13217 (n7124, n6814, n7123);
  not g13218 (n_6343, n7124);
  and g13219 (n7125, n6814, n_6343);
  and g13220 (n7126, n7123, n_6343);
  not g13221 (n_6344, n7125);
  not g13222 (n_6345, n7126);
  and g13223 (n7127, n_6344, n_6345);
  not g13224 (n_6346, n6932);
  not g13225 (n_6347, n7127);
  and g13226 (n7128, n_6346, n_6347);
  not g13227 (n_6348, n7128);
  and g13228 (n7129, n_6346, n_6348);
  and g13229 (n7130, n_6347, n_6348);
  not g13230 (n_6349, n7129);
  not g13231 (n_6350, n7130);
  and g13232 (n7131, n_6349, n_6350);
  not g13233 (n_6351, n7131);
  and g13234 (n7132, n7118, n_6351);
  not g13235 (n_6352, n7132);
  and g13236 (n7133, n7118, n_6352);
  and g13237 (n7134, n_6351, n_6352);
  not g13238 (n_6353, n7133);
  not g13239 (n_6354, n7134);
  and g13240 (n7135, n_6353, n_6354);
  and g13241 (n7136, n_6200, n_6244);
  not g13242 (n_6355, n7135);
  not g13243 (n_6356, n7136);
  and g13244 (n7137, n_6355, n_6356);
  not g13245 (n_6357, n7137);
  and g13246 (n7138, n_6355, n_6357);
  and g13247 (n7139, n_6356, n_6357);
  not g13248 (n_6358, n7138);
  not g13249 (n_6359, n7139);
  and g13250 (n7140, n_6358, n_6359);
  and g13251 (n7141, n_6054, n_6062);
  and g13252 (n7142, n6989, n7141);
  not g13253 (n_6360, n6989);
  not g13254 (n_6361, n7141);
  and g13255 (n7143, n_6360, n_6361);
  not g13256 (n_6362, n7142);
  not g13257 (n_6363, n7143);
  and g13258 (n7144, n_6362, n_6363);
  and g13259 (n7145, \a[18] , \a[37] );
  and g13260 (n7146, \a[19] , \a[36] );
  not g13261 (n_6364, n7145);
  not g13262 (n_6365, n7146);
  and g13263 (n7147, n_6364, n_6365);
  and g13264 (n7148, n1149, n3687);
  not g13265 (n_6366, n7148);
  not g13268 (n_6367, n7147);
  not g13270 (n_6368, n7151);
  and g13271 (n7152, \a[50] , n_6368);
  and g13272 (n7153, \a[5] , n7152);
  and g13273 (n7154, n_6366, n_6368);
  and g13274 (n7155, n_6367, n7154);
  not g13275 (n_6369, n7153);
  not g13276 (n_6370, n7155);
  and g13277 (n7156, n_6369, n_6370);
  not g13278 (n_6371, n7156);
  and g13279 (n7157, n7144, n_6371);
  not g13280 (n_6372, n7157);
  and g13281 (n7158, n7144, n_6372);
  and g13282 (n7159, n_6371, n_6372);
  not g13283 (n_6373, n7158);
  not g13284 (n_6374, n7159);
  and g13285 (n7160, n_6373, n_6374);
  and g13286 (n7161, n6972, n7004);
  not g13287 (n_6375, n6972);
  not g13288 (n_6376, n7004);
  and g13289 (n7162, n_6375, n_6376);
  not g13290 (n_6377, n7161);
  not g13291 (n_6378, n7162);
  and g13292 (n7163, n_6377, n_6378);
  not g13293 (n_6379, n7163);
  and g13294 (n7164, n6920, n_6379);
  not g13295 (n_6380, n6920);
  and g13296 (n7165, n_6380, n7163);
  not g13297 (n_6381, n7164);
  not g13298 (n_6382, n7165);
  and g13299 (n7166, n_6381, n_6382);
  and g13300 (n7167, n_6090, n_6091);
  not g13301 (n_6383, n7167);
  and g13302 (n7168, n_6087, n_6383);
  not g13303 (n_6384, n7168);
  and g13304 (n7169, n7166, n_6384);
  not g13305 (n_6385, n7166);
  and g13306 (n7170, n_6385, n7168);
  not g13307 (n_6386, n7169);
  not g13308 (n_6387, n7170);
  and g13309 (n7171, n_6386, n_6387);
  not g13310 (n_6388, n7160);
  and g13311 (n7172, n_6388, n7171);
  not g13312 (n_6389, n7172);
  and g13313 (n7173, n_6388, n_6389);
  and g13314 (n7174, n7171, n_6389);
  not g13315 (n_6390, n7173);
  not g13316 (n_6391, n7174);
  and g13317 (n7175, n_6390, n_6391);
  not g13318 (n_6392, n7140);
  not g13319 (n_6393, n7175);
  and g13320 (n7176, n_6392, n_6393);
  not g13321 (n_6394, n7176);
  and g13322 (n7177, n_6392, n_6394);
  and g13323 (n7178, n_6393, n_6394);
  not g13324 (n_6395, n7177);
  not g13325 (n_6396, n7178);
  and g13326 (n7179, n_6395, n_6396);
  and g13327 (n7180, n_6052, n_6105);
  and g13328 (n7181, n7179, n7180);
  not g13329 (n_6397, n7179);
  not g13330 (n_6398, n7180);
  and g13331 (n7182, n_6397, n_6398);
  not g13332 (n_6399, n7181);
  not g13333 (n_6400, n7182);
  and g13334 (n7183, n_6399, n_6400);
  and g13335 (n7184, n818, n4639);
  and g13336 (n7185, n723, n5713);
  and g13337 (n7186, \a[13] , \a[45] );
  and g13338 (n7187, n6451, n7186);
  not g13339 (n_6401, n7185);
  not g13340 (n_6402, n7187);
  and g13341 (n7188, n_6401, n_6402);
  not g13342 (n_6403, n7184);
  not g13343 (n_6404, n7188);
  and g13344 (n7189, n_6403, n_6404);
  not g13345 (n_6405, n7189);
  and g13346 (n7190, n_6403, n_6405);
  and g13347 (n7191, \a[11] , \a[44] );
  not g13348 (n_6406, n5949);
  not g13349 (n_6407, n7191);
  and g13350 (n7192, n_6406, n_6407);
  not g13351 (n_6408, n7192);
  and g13352 (n7193, n7190, n_6408);
  and g13353 (n7194, \a[45] , n_6405);
  and g13354 (n7195, \a[10] , n7194);
  not g13355 (n_6409, n7193);
  not g13356 (n_6410, n7195);
  and g13357 (n7196, n_6409, n_6410);
  and g13358 (n7197, \a[26] , \a[29] );
  not g13359 (n_6411, n2331);
  not g13360 (n_6412, n7197);
  and g13361 (n7198, n_6411, n_6412);
  and g13362 (n7199, n2331, n7197);
  not g13363 (n_6413, n7199);
  not g13366 (n_6414, n7198);
  not g13368 (n_6415, n7202);
  and g13369 (n7203, \a[43] , n_6415);
  and g13370 (n7204, \a[12] , n7203);
  and g13371 (n7205, n_6413, n_6415);
  and g13372 (n7206, n_6414, n7205);
  not g13373 (n_6416, n7204);
  not g13374 (n_6417, n7206);
  and g13375 (n7207, n_6416, n_6417);
  not g13376 (n_6418, n7196);
  not g13377 (n_6419, n7207);
  and g13378 (n7208, n_6418, n_6419);
  not g13379 (n_6420, n7208);
  and g13380 (n7209, n_6418, n_6420);
  and g13381 (n7210, n_6419, n_6420);
  not g13382 (n_6421, n7209);
  not g13383 (n_6422, n7210);
  and g13384 (n7211, n_6421, n_6422);
  and g13385 (n7212, \a[7] , \a[48] );
  and g13386 (n7213, \a[8] , \a[47] );
  not g13387 (n_6423, n7212);
  not g13388 (n_6424, n7213);
  and g13389 (n7214, n_6423, n_6424);
  and g13390 (n7215, n380, n6252);
  not g13391 (n_6425, n7215);
  not g13394 (n_6426, n7214);
  not g13396 (n_6427, n7218);
  and g13397 (n7219, \a[39] , n_6427);
  and g13398 (n7220, \a[16] , n7219);
  and g13399 (n7221, n_6425, n_6427);
  and g13400 (n7222, n_6426, n7221);
  not g13401 (n_6428, n7220);
  not g13402 (n_6429, n7222);
  and g13403 (n7223, n_6428, n_6429);
  not g13404 (n_6430, n7211);
  not g13405 (n_6431, n7223);
  and g13406 (n7224, n_6430, n_6431);
  not g13407 (n_6432, n7224);
  and g13408 (n7225, n_6430, n_6432);
  and g13409 (n7226, n_6431, n_6432);
  not g13410 (n_6433, n7225);
  not g13411 (n_6434, n7226);
  and g13412 (n7227, n_6433, n_6434);
  and g13413 (n7228, n_6116, n_6120);
  and g13414 (n7229, n7227, n7228);
  not g13415 (n_6435, n7227);
  not g13416 (n_6436, n7228);
  and g13417 (n7230, n_6435, n_6436);
  not g13418 (n_6437, n7229);
  not g13419 (n_6438, n7230);
  and g13420 (n7231, n_6437, n_6438);
  and g13421 (n7232, \a[51] , \a[53] );
  and g13422 (n7233, n252, n7232);
  and g13423 (n7234, \a[51] , n212);
  and g13424 (n7235, \a[53] , n196);
  not g13425 (n_6439, n7234);
  not g13426 (n_6440, n7235);
  and g13427 (n7236, n_6439, n_6440);
  not g13428 (n_6442, n7233);
  and g13429 (n7237, \a[55] , n_6442);
  not g13430 (n_6443, n7236);
  and g13431 (n7238, n_6443, n7237);
  not g13432 (n_6444, n7238);
  and g13433 (n7239, n_6442, n_6444);
  and g13434 (n7240, \a[2] , \a[53] );
  and g13435 (n7241, \a[4] , \a[51] );
  not g13436 (n_6445, n7240);
  not g13437 (n_6446, n7241);
  and g13438 (n7242, n_6445, n_6446);
  not g13439 (n_6447, n7242);
  and g13440 (n7243, n7239, n_6447);
  and g13441 (n7244, \a[55] , n_6444);
  and g13442 (n7245, \a[0] , n7244);
  not g13443 (n_6448, n7243);
  not g13444 (n_6449, n7245);
  and g13445 (n7246, n_6448, n_6449);
  and g13446 (n7247, n1574, n4150);
  and g13447 (n7248, n1693, n2972);
  and g13448 (n7249, n1494, n3319);
  not g13449 (n_6450, n7248);
  not g13450 (n_6451, n7249);
  and g13451 (n7250, n_6450, n_6451);
  not g13452 (n_6452, n7247);
  not g13453 (n_6453, n7250);
  and g13454 (n7251, n_6452, n_6453);
  not g13455 (n_6454, n7251);
  and g13456 (n7252, \a[35] , n_6454);
  and g13457 (n7253, \a[20] , n7252);
  and g13458 (n7254, n_6452, n_6454);
  and g13459 (n7255, \a[21] , \a[34] );
  not g13460 (n_6455, n2595);
  not g13461 (n_6456, n7255);
  and g13462 (n7256, n_6455, n_6456);
  not g13463 (n_6457, n7256);
  and g13464 (n7257, n7254, n_6457);
  not g13465 (n_6458, n7253);
  not g13466 (n_6459, n7257);
  and g13467 (n7258, n_6458, n_6459);
  not g13468 (n_6460, n7246);
  not g13469 (n_6461, n7258);
  and g13470 (n7259, n_6460, n_6461);
  not g13471 (n_6462, n7259);
  and g13472 (n7260, n_6460, n_6462);
  and g13473 (n7261, n_6461, n_6462);
  not g13474 (n_6463, n7260);
  not g13475 (n_6464, n7261);
  and g13476 (n7262, n_6463, n_6464);
  and g13477 (n7263, \a[23] , \a[32] );
  and g13478 (n7264, n1904, n2865);
  and g13479 (n7265, n1547, n2488);
  and g13480 (n7266, n1666, n3812);
  not g13481 (n_6465, n7265);
  not g13482 (n_6466, n7266);
  and g13483 (n7267, n_6465, n_6466);
  not g13484 (n_6467, n7264);
  not g13485 (n_6468, n7267);
  and g13486 (n7268, n_6467, n_6468);
  not g13487 (n_6469, n7268);
  and g13488 (n7269, n7263, n_6469);
  and g13489 (n7270, n_6467, n_6469);
  and g13490 (n7271, \a[24] , \a[31] );
  and g13491 (n7272, \a[25] , \a[30] );
  not g13492 (n_6470, n7271);
  not g13493 (n_6471, n7272);
  and g13494 (n7273, n_6470, n_6471);
  not g13495 (n_6472, n7273);
  and g13496 (n7274, n7270, n_6472);
  not g13497 (n_6473, n7269);
  not g13498 (n_6474, n7274);
  and g13499 (n7275, n_6473, n_6474);
  not g13500 (n_6475, n7262);
  not g13501 (n_6476, n7275);
  and g13502 (n7276, n_6475, n_6476);
  not g13503 (n_6477, n7276);
  and g13504 (n7277, n_6475, n_6477);
  and g13505 (n7278, n_6476, n_6477);
  not g13506 (n_6478, n7277);
  not g13507 (n_6479, n7278);
  and g13508 (n7279, n_6478, n_6479);
  not g13509 (n_6480, n7279);
  and g13510 (n7280, n7231, n_6480);
  not g13511 (n_6481, n7231);
  and g13512 (n7281, n_6481, n7279);
  and g13513 (n7282, n_6096, n_6101);
  and g13514 (n7283, n6828, n6843);
  not g13515 (n_6482, n6828);
  not g13516 (n_6483, n6843);
  and g13517 (n7284, n_6482, n_6483);
  not g13518 (n_6484, n7283);
  not g13519 (n_6485, n7284);
  and g13520 (n7285, n_6484, n_6485);
  not g13521 (n_6486, n7285);
  and g13522 (n7286, n6954, n_6486);
  not g13523 (n_6487, n6954);
  and g13524 (n7287, n_6487, n7285);
  not g13525 (n_6488, n7286);
  not g13526 (n_6489, n7287);
  and g13527 (n7288, n_6488, n_6489);
  and g13528 (n7289, n_6179, n_6194);
  and g13529 (n7290, n_6223, n_6238);
  and g13530 (n7291, n7289, n7290);
  not g13531 (n_6490, n7289);
  not g13532 (n_6491, n7290);
  and g13533 (n7292, n_6490, n_6491);
  not g13534 (n_6492, n7291);
  not g13535 (n_6493, n7292);
  and g13536 (n7293, n_6492, n_6493);
  and g13537 (n7294, n7288, n7293);
  not g13538 (n_6494, n7288);
  not g13539 (n_6495, n7293);
  and g13540 (n7295, n_6494, n_6495);
  not g13541 (n_6496, n7294);
  not g13542 (n_6497, n7295);
  and g13543 (n7296, n_6496, n_6497);
  not g13544 (n_6498, n7282);
  and g13545 (n7297, n_6498, n7296);
  not g13546 (n_6499, n7296);
  and g13547 (n7298, n7282, n_6499);
  not g13548 (n_6500, n7297);
  not g13549 (n_6501, n7298);
  and g13550 (n7299, n_6500, n_6501);
  not g13551 (n_6502, n7281);
  and g13552 (n7300, n_6502, n7299);
  not g13553 (n_6503, n7280);
  and g13554 (n7301, n_6503, n7300);
  not g13555 (n_6504, n7301);
  and g13556 (n7302, n7299, n_6504);
  and g13557 (n7303, n_6502, n_6504);
  and g13558 (n7304, n_6503, n7303);
  not g13559 (n_6505, n7302);
  not g13560 (n_6506, n7304);
  and g13561 (n7305, n_6505, n_6506);
  not g13562 (n_6507, n7183);
  and g13563 (n7306, n_6507, n7305);
  not g13564 (n_6508, n7305);
  and g13565 (n7307, n7183, n_6508);
  not g13566 (n_6509, n7306);
  not g13567 (n_6510, n7307);
  and g13568 (n7308, n_6509, n_6510);
  not g13569 (n_6511, n7113);
  and g13570 (n7309, n_6511, n7308);
  not g13571 (n_6512, n7308);
  and g13572 (n7310, n7113, n_6512);
  not g13573 (n_6513, n7309);
  not g13574 (n_6514, n7310);
  and g13575 (n7311, n_6513, n_6514);
  not g13576 (n_6515, n7055);
  and g13577 (n7312, n_6515, n7311);
  not g13578 (n_6516, n7311);
  and g13579 (n7313, n7055, n_6516);
  not g13580 (n_6517, n7312);
  not g13581 (n_6518, n7313);
  and g13582 (n7314, n_6517, n_6518);
  and g13583 (n7315, n_6280, n_6283);
  not g13584 (n_6519, n7315);
  and g13585 (n7316, n_6279, n_6519);
  not g13586 (n_6520, n7314);
  and g13587 (n7317, n_6520, n7316);
  not g13588 (n_6521, n7316);
  and g13589 (n7318, n7314, n_6521);
  not g13590 (n_6522, n7317);
  not g13591 (n_6523, n7318);
  and g13592 (\asquared[56] , n_6522, n_6523);
  and g13593 (n7320, n_6332, n_6513);
  and g13594 (n7321, \a[7] , \a[49] );
  and g13595 (n7322, \a[17] , \a[39] );
  not g13596 (n_6524, n7321);
  not g13597 (n_6525, n7322);
  and g13598 (n7323, n_6524, n_6525);
  and g13599 (n7324, n335, n6325);
  and g13600 (n7325, \a[17] , \a[50] );
  and g13601 (n7326, n4746, n7325);
  not g13602 (n_6526, n7324);
  not g13603 (n_6527, n7326);
  and g13604 (n7327, n_6526, n_6527);
  and g13605 (n7328, n7321, n7322);
  not g13606 (n_6528, n7327);
  not g13607 (n_6529, n7328);
  and g13608 (n7329, n_6528, n_6529);
  not g13609 (n_6530, n7329);
  and g13610 (n7330, n_6529, n_6530);
  not g13611 (n_6531, n7323);
  and g13612 (n7331, n_6531, n7330);
  and g13613 (n7332, \a[50] , n_6530);
  and g13614 (n7333, \a[6] , n7332);
  not g13615 (n_6532, n7331);
  not g13616 (n_6533, n7333);
  and g13617 (n7334, n_6532, n_6533);
  and g13618 (n7335, n748, n5296);
  and g13619 (n7336, n818, n4811);
  and g13620 (n7337, n602, n5713);
  not g13621 (n_6534, n7336);
  not g13622 (n_6535, n7337);
  and g13623 (n7338, n_6534, n_6535);
  not g13624 (n_6536, n7335);
  not g13625 (n_6537, n7338);
  and g13626 (n7339, n_6536, n_6537);
  not g13627 (n_6538, n7339);
  and g13628 (n7340, \a[45] , n_6538);
  and g13629 (n7341, \a[11] , n7340);
  and g13630 (n7342, \a[12] , \a[44] );
  not g13631 (n_6539, n6165);
  not g13632 (n_6540, n7342);
  and g13633 (n7343, n_6539, n_6540);
  and g13634 (n7344, n_6536, n_6538);
  not g13635 (n_6541, n7343);
  and g13636 (n7345, n_6541, n7344);
  not g13637 (n_6542, n7341);
  not g13638 (n_6543, n7345);
  and g13639 (n7346, n_6542, n_6543);
  not g13640 (n_6544, n7334);
  not g13641 (n_6545, n7346);
  and g13642 (n7347, n_6544, n_6545);
  not g13643 (n_6546, n7347);
  and g13644 (n7348, n_6544, n_6546);
  and g13645 (n7349, n_6545, n_6546);
  not g13646 (n_6547, n7348);
  not g13647 (n_6548, n7349);
  and g13648 (n7350, n_6547, n_6548);
  and g13649 (n7351, \a[15] , \a[48] );
  and g13650 (n7352, n5620, n7351);
  and g13651 (n7353, \a[40] , \a[48] );
  and g13652 (n7354, n1509, n7353);
  and g13653 (n7355, n891, n5413);
  not g13654 (n_6549, n7354);
  not g13655 (n_6550, n7355);
  and g13656 (n7356, n_6549, n_6550);
  not g13657 (n_6551, n7352);
  not g13658 (n_6552, n7356);
  and g13659 (n7357, n_6551, n_6552);
  not g13660 (n_6553, n7357);
  and g13661 (n7358, n4169, n_6553);
  and g13662 (n7359, n_6551, n_6553);
  and g13663 (n7360, \a[8] , \a[48] );
  and g13664 (n7361, \a[15] , \a[41] );
  not g13665 (n_6554, n7360);
  not g13666 (n_6555, n7361);
  and g13667 (n7362, n_6554, n_6555);
  not g13668 (n_6556, n7362);
  and g13669 (n7363, n7359, n_6556);
  not g13670 (n_6557, n7358);
  not g13671 (n_6558, n7363);
  and g13672 (n7364, n_6557, n_6558);
  not g13673 (n_6559, n7350);
  not g13674 (n_6560, n7364);
  and g13675 (n7365, n_6559, n_6560);
  not g13676 (n_6561, n7365);
  and g13677 (n7366, n_6559, n_6561);
  and g13678 (n7367, n_6560, n_6561);
  not g13679 (n_6562, n7366);
  not g13680 (n_6563, n7367);
  and g13681 (n7368, n_6562, n_6563);
  and g13682 (n7369, n1919, n4150);
  and g13683 (n7370, n1693, n4595);
  and g13684 (n7371, \a[33] , \a[36] );
  and g13685 (n7372, n4423, n7371);
  not g13686 (n_6564, n7370);
  not g13687 (n_6565, n7372);
  and g13688 (n7373, n_6564, n_6565);
  not g13689 (n_6566, n7369);
  not g13690 (n_6567, n7373);
  and g13691 (n7374, n_6566, n_6567);
  not g13692 (n_6568, n7374);
  and g13693 (n7375, n_6566, n_6568);
  and g13694 (n7376, \a[22] , \a[34] );
  and g13695 (n7377, \a[23] , \a[33] );
  not g13696 (n_6569, n7376);
  not g13697 (n_6570, n7377);
  and g13698 (n7378, n_6569, n_6570);
  not g13699 (n_6571, n7378);
  and g13700 (n7379, n7375, n_6571);
  and g13701 (n7380, \a[36] , n_6568);
  and g13702 (n7381, \a[20] , n7380);
  not g13703 (n_6572, n7379);
  not g13704 (n_6573, n7381);
  and g13705 (n7382, n_6572, n_6573);
  and g13706 (n7383, n2463, n2865);
  and g13707 (n7384, n2301, n2488);
  and g13708 (n7385, n1904, n3812);
  not g13709 (n_6574, n7384);
  not g13710 (n_6575, n7385);
  and g13711 (n7386, n_6574, n_6575);
  not g13712 (n_6576, n7383);
  not g13713 (n_6577, n7386);
  and g13714 (n7387, n_6576, n_6577);
  not g13715 (n_6578, n7387);
  and g13716 (n7388, \a[32] , n_6578);
  and g13717 (n7389, \a[24] , n7388);
  and g13718 (n7390, n_6576, n_6578);
  and g13719 (n7391, \a[25] , \a[31] );
  and g13720 (n7392, \a[26] , \a[30] );
  not g13721 (n_6579, n7391);
  not g13722 (n_6580, n7392);
  and g13723 (n7393, n_6579, n_6580);
  not g13724 (n_6581, n7393);
  and g13725 (n7394, n7390, n_6581);
  not g13726 (n_6582, n7389);
  not g13727 (n_6583, n7394);
  and g13728 (n7395, n_6582, n_6583);
  not g13729 (n_6584, n7382);
  not g13730 (n_6585, n7395);
  and g13731 (n7396, n_6584, n_6585);
  not g13732 (n_6586, n7396);
  and g13733 (n7397, n_6584, n_6586);
  and g13734 (n7398, n_6585, n_6586);
  not g13735 (n_6587, n7397);
  not g13736 (n_6588, n7398);
  and g13737 (n7399, n_6587, n_6588);
  and g13738 (n7400, \a[14] , \a[46] );
  and g13739 (n7401, n6451, n7400);
  and g13740 (n7402, n484, n5666);
  and g13741 (n7403, \a[14] , \a[47] );
  and g13742 (n7404, n6180, n7403);
  not g13743 (n_6589, n7402);
  not g13744 (n_6590, n7404);
  and g13745 (n7405, n_6589, n_6590);
  not g13746 (n_6591, n7401);
  not g13747 (n_6592, n7405);
  and g13748 (n7406, n_6591, n_6592);
  not g13749 (n_6593, n7406);
  and g13750 (n7407, \a[47] , n_6593);
  and g13751 (n7408, \a[9] , n7407);
  and g13752 (n7409, n_6591, n_6593);
  and g13753 (n7410, \a[10] , \a[46] );
  not g13754 (n_6594, n5346);
  not g13755 (n_6595, n7410);
  and g13756 (n7411, n_6594, n_6595);
  not g13757 (n_6596, n7411);
  and g13758 (n7412, n7409, n_6596);
  not g13759 (n_6597, n7408);
  not g13760 (n_6598, n7412);
  and g13761 (n7413, n_6597, n_6598);
  not g13762 (n_6599, n7399);
  not g13763 (n_6600, n7413);
  and g13764 (n7414, n_6599, n_6600);
  not g13765 (n_6601, n7414);
  and g13766 (n7415, n_6599, n_6601);
  and g13767 (n7416, n_6600, n_6601);
  not g13768 (n_6602, n7415);
  not g13769 (n_6603, n7416);
  and g13770 (n7417, n_6602, n_6603);
  not g13771 (n_6604, n7368);
  and g13772 (n7418, n_6604, n7417);
  not g13773 (n_6605, n7417);
  and g13774 (n7419, n7368, n_6605);
  not g13775 (n_6606, n7418);
  not g13776 (n_6607, n7419);
  and g13777 (n7420, n_6606, n_6607);
  and g13778 (n7421, \a[54] , \a[56] );
  and g13779 (n7422, n196, n7421);
  and g13780 (n7423, \a[0] , \a[56] );
  and g13781 (n7424, \a[2] , \a[54] );
  not g13782 (n_6609, n7423);
  not g13783 (n_6610, n7424);
  and g13784 (n7425, n_6609, n_6610);
  not g13785 (n_6611, n7422);
  not g13786 (n_6612, n7425);
  and g13787 (n7426, n_6611, n_6612);
  and g13788 (n7427, n7120, n7426);
  not g13789 (n_6613, n7426);
  and g13790 (n7428, n_6341, n_6613);
  not g13791 (n_6614, n7427);
  not g13792 (n_6615, n7428);
  and g13793 (n7429, n_6614, n_6615);
  not g13794 (n_6616, n7221);
  and g13795 (n7430, n_6616, n7429);
  not g13796 (n_6617, n7429);
  and g13797 (n7431, n7221, n_6617);
  not g13798 (n_6618, n7430);
  not g13799 (n_6619, n7431);
  and g13800 (n7432, n_6618, n_6619);
  and g13801 (n7433, \a[52] , \a[53] );
  and g13802 (n7434, n209, n7433);
  and g13803 (n7435, \a[37] , \a[53] );
  and g13804 (n7436, n1273, n7435);
  not g13805 (n_6620, n7434);
  not g13806 (n_6621, n7436);
  and g13807 (n7437, n_6620, n_6621);
  and g13808 (n7438, \a[4] , \a[52] );
  and g13809 (n7439, \a[19] , \a[37] );
  and g13810 (n7440, n7438, n7439);
  not g13811 (n_6622, n7437);
  not g13812 (n_6623, n7440);
  and g13813 (n7441, n_6622, n_6623);
  not g13814 (n_6624, n7441);
  and g13815 (n7442, \a[53] , n_6624);
  and g13816 (n7443, \a[3] , n7442);
  and g13817 (n7444, n_6623, n_6624);
  not g13818 (n_6625, n7438);
  not g13819 (n_6626, n7439);
  and g13820 (n7445, n_6625, n_6626);
  not g13821 (n_6627, n7445);
  and g13822 (n7446, n7444, n_6627);
  not g13823 (n_6628, n7443);
  not g13824 (n_6629, n7446);
  and g13825 (n7447, n_6628, n_6629);
  not g13826 (n_6630, n7447);
  and g13827 (n7448, n7432, n_6630);
  not g13828 (n_6631, n7448);
  and g13829 (n7449, n7432, n_6631);
  and g13830 (n7450, n_6630, n_6631);
  not g13831 (n_6632, n7449);
  not g13832 (n_6633, n7450);
  and g13833 (n7451, n_6632, n_6633);
  and g13834 (n7452, n7420, n7451);
  not g13835 (n_6634, n7420);
  not g13836 (n_6635, n7451);
  and g13837 (n7453, n_6634, n_6635);
  not g13838 (n_6636, n7452);
  not g13839 (n_6637, n7453);
  and g13840 (n7454, n_6636, n_6637);
  and g13841 (n7455, n_6315, n_6319);
  and g13842 (n7456, n7254, n7270);
  not g13843 (n_6638, n7254);
  not g13844 (n_6639, n7270);
  and g13845 (n7457, n_6638, n_6639);
  not g13846 (n_6640, n7456);
  not g13847 (n_6641, n7457);
  and g13848 (n7458, n_6640, n_6641);
  not g13849 (n_6642, n7458);
  and g13850 (n7459, n7068, n_6642);
  not g13851 (n_6643, n7068);
  and g13852 (n7460, n_6643, n7458);
  not g13853 (n_6644, n7459);
  not g13854 (n_6645, n7460);
  and g13855 (n7461, n_6644, n_6645);
  and g13856 (n7462, n_6420, n_6432);
  and g13857 (n7463, \a[1] , \a[55] );
  not g13858 (n_6646, n2041);
  not g13859 (n_6647, n7463);
  and g13860 (n7464, n_6646, n_6647);
  and g13861 (n7465, n2041, n7463);
  not g13862 (n_6648, n7205);
  not g13863 (n_6649, n7465);
  and g13864 (n7466, n_6648, n_6649);
  not g13865 (n_6650, n7464);
  and g13866 (n7467, n_6650, n7466);
  not g13867 (n_6651, n7467);
  and g13868 (n7468, n_6648, n_6651);
  and g13869 (n7469, n_6649, n_6651);
  and g13870 (n7470, n_6650, n7469);
  not g13871 (n_6652, n7468);
  not g13872 (n_6653, n7470);
  and g13873 (n7471, n_6652, n_6653);
  not g13874 (n_6654, n7190);
  not g13875 (n_6655, n7471);
  and g13876 (n7472, n_6654, n_6655);
  and g13877 (n7473, n7190, n_6653);
  and g13878 (n7474, n_6652, n7473);
  not g13879 (n_6656, n7472);
  not g13880 (n_6657, n7474);
  and g13881 (n7475, n_6656, n_6657);
  not g13882 (n_6658, n7462);
  and g13883 (n7476, n_6658, n7475);
  not g13884 (n_6659, n7475);
  and g13885 (n7477, n7462, n_6659);
  not g13886 (n_6660, n7476);
  not g13887 (n_6661, n7477);
  and g13888 (n7478, n_6660, n_6661);
  and g13889 (n7479, n7461, n7478);
  not g13890 (n_6662, n7461);
  not g13891 (n_6663, n7478);
  and g13892 (n7480, n_6662, n_6663);
  not g13893 (n_6664, n7479);
  not g13894 (n_6665, n7480);
  and g13895 (n7481, n_6664, n_6665);
  not g13896 (n_6666, n7455);
  and g13897 (n7482, n_6666, n7481);
  not g13898 (n_6667, n7482);
  and g13899 (n7483, n_6666, n_6667);
  and g13900 (n7484, n7481, n_6667);
  not g13901 (n_6668, n7483);
  not g13902 (n_6669, n7484);
  and g13903 (n7485, n_6668, n_6669);
  not g13904 (n_6670, n7485);
  and g13905 (n7486, n7454, n_6670);
  not g13906 (n_6671, n7486);
  and g13907 (n7487, n7454, n_6671);
  and g13908 (n7488, n_6670, n_6671);
  not g13909 (n_6672, n7487);
  not g13910 (n_6673, n7488);
  and g13911 (n7489, n_6672, n_6673);
  and g13912 (n7490, n_6322, n_6327);
  and g13913 (n7491, n7154, n7239);
  not g13914 (n_6674, n7154);
  not g13915 (n_6675, n7239);
  and g13916 (n7492, n_6674, n_6675);
  not g13917 (n_6676, n7491);
  not g13918 (n_6677, n7492);
  and g13919 (n7493, n_6676, n_6677);
  not g13920 (n_6678, n7493);
  and g13921 (n7494, n7084, n_6678);
  not g13922 (n_6679, n7084);
  and g13923 (n7495, n_6679, n7493);
  not g13924 (n_6680, n7494);
  not g13925 (n_6681, n7495);
  and g13926 (n7496, n_6680, n_6681);
  and g13927 (n7497, n_6306, n_6312);
  not g13928 (n_6682, n7496);
  and g13929 (n7498, n_6682, n7497);
  not g13930 (n_6683, n7497);
  and g13931 (n7499, n7496, n_6683);
  not g13932 (n_6684, n7498);
  not g13933 (n_6685, n7499);
  and g13934 (n7500, n_6684, n_6685);
  and g13935 (n7501, n_6338, n_6352);
  not g13936 (n_6686, n7500);
  and g13937 (n7502, n_6686, n7501);
  not g13938 (n_6687, n7501);
  and g13939 (n7503, n7500, n_6687);
  not g13940 (n_6688, n7502);
  not g13941 (n_6689, n7503);
  and g13942 (n7504, n_6688, n_6689);
  and g13943 (n7505, n_6485, n_6489);
  and g13944 (n7506, n_6363, n_6372);
  and g13945 (n7507, n7505, n7506);
  not g13946 (n_6690, n7505);
  not g13947 (n_6691, n7506);
  and g13948 (n7508, n_6690, n_6691);
  not g13949 (n_6692, n7507);
  not g13950 (n_6693, n7508);
  and g13951 (n7509, n_6692, n_6693);
  and g13952 (n7510, n_6462, n_6477);
  not g13953 (n_6694, n7509);
  and g13954 (n7511, n_6694, n7510);
  not g13955 (n_6695, n7510);
  and g13956 (n7512, n7509, n_6695);
  not g13957 (n_6696, n7511);
  not g13958 (n_6697, n7512);
  and g13959 (n7513, n_6696, n_6697);
  and g13960 (n7514, n_6438, n_6503);
  not g13961 (n_6698, n7514);
  and g13962 (n7515, n7513, n_6698);
  not g13963 (n_6699, n7515);
  and g13964 (n7516, n7513, n_6699);
  and g13965 (n7517, n_6698, n_6699);
  not g13966 (n_6700, n7516);
  not g13967 (n_6701, n7517);
  and g13968 (n7518, n_6700, n_6701);
  not g13969 (n_6702, n7518);
  and g13970 (n7519, n7504, n_6702);
  not g13971 (n_6703, n7504);
  and g13972 (n7520, n_6703, n_6701);
  and g13973 (n7521, n_6700, n7520);
  not g13974 (n_6704, n7519);
  not g13975 (n_6705, n7521);
  and g13976 (n7522, n_6704, n_6705);
  not g13977 (n_6706, n7490);
  and g13978 (n7523, n_6706, n7522);
  not g13979 (n_6707, n7523);
  and g13980 (n7524, n_6706, n_6707);
  and g13981 (n7525, n7522, n_6707);
  not g13982 (n_6708, n7524);
  not g13983 (n_6709, n7525);
  and g13984 (n7526, n_6708, n_6709);
  not g13985 (n_6710, n7489);
  not g13986 (n_6711, n7526);
  and g13987 (n7527, n_6710, n_6711);
  not g13988 (n_6712, n7527);
  and g13989 (n7528, n_6710, n_6712);
  and g13990 (n7529, n_6711, n_6712);
  not g13991 (n_6713, n7528);
  not g13992 (n_6714, n7529);
  and g13993 (n7530, n_6713, n_6714);
  and g13994 (n7531, n_6386, n_6389);
  and g13995 (n7532, n_6343, n_6348);
  and g13996 (n7533, \a[5] , \a[51] );
  and g13997 (n7534, \a[18] , \a[38] );
  not g13998 (n_6715, n7533);
  not g13999 (n_6716, n7534);
  and g14000 (n7535, n_6715, n_6716);
  and g14001 (n7536, \a[38] , \a[51] );
  and g14002 (n7537, n1340, n7536);
  not g14003 (n_6717, n7537);
  not g14006 (n_6718, n7535);
  not g14008 (n_6719, n7540);
  and g14009 (n7541, \a[35] , n_6719);
  and g14010 (n7542, \a[21] , n7541);
  and g14011 (n7543, n_6717, n_6719);
  and g14012 (n7544, n_6718, n7543);
  not g14013 (n_6720, n7542);
  not g14014 (n_6721, n7544);
  and g14015 (n7545, n_6720, n_6721);
  not g14016 (n_6722, n7532);
  not g14017 (n_6723, n7545);
  and g14018 (n7546, n_6722, n_6723);
  not g14019 (n_6724, n7546);
  and g14020 (n7547, n_6722, n_6724);
  and g14021 (n7548, n_6723, n_6724);
  not g14022 (n_6725, n7547);
  not g14023 (n_6726, n7548);
  and g14024 (n7549, n_6725, n_6726);
  and g14025 (n7550, n_6378, n_6382);
  and g14026 (n7551, n7549, n7550);
  not g14027 (n_6727, n7549);
  not g14028 (n_6728, n7550);
  and g14029 (n7552, n_6727, n_6728);
  not g14030 (n_6729, n7551);
  not g14031 (n_6730, n7552);
  and g14032 (n7553, n_6729, n_6730);
  and g14033 (n7554, n_6493, n_6496);
  not g14034 (n_6731, n7554);
  and g14035 (n7555, n7553, n_6731);
  not g14036 (n_6732, n7553);
  and g14037 (n7556, n_6732, n7554);
  not g14038 (n_6733, n7555);
  not g14039 (n_6734, n7556);
  and g14040 (n7557, n_6733, n_6734);
  not g14041 (n_6735, n7557);
  and g14042 (n7558, n7531, n_6735);
  not g14043 (n_6736, n7531);
  and g14044 (n7559, n_6736, n7557);
  not g14045 (n_6737, n7558);
  not g14046 (n_6738, n7559);
  and g14047 (n7560, n_6737, n_6738);
  and g14048 (n7561, n_6357, n_6394);
  not g14049 (n_6739, n7560);
  and g14050 (n7562, n_6739, n7561);
  not g14051 (n_6740, n7561);
  and g14052 (n7563, n7560, n_6740);
  not g14053 (n_6741, n7562);
  not g14054 (n_6742, n7563);
  and g14055 (n7564, n_6741, n_6742);
  and g14056 (n7565, n_6500, n_6504);
  not g14057 (n_6743, n7564);
  and g14058 (n7566, n_6743, n7565);
  not g14059 (n_6744, n7565);
  and g14060 (n7567, n7564, n_6744);
  not g14061 (n_6745, n7566);
  not g14062 (n_6746, n7567);
  and g14063 (n7568, n_6745, n_6746);
  and g14064 (n7569, n_6400, n_6510);
  not g14065 (n_6747, n7569);
  and g14066 (n7570, n7568, n_6747);
  not g14067 (n_6748, n7570);
  and g14068 (n7571, n7568, n_6748);
  and g14069 (n7572, n_6747, n_6748);
  not g14070 (n_6749, n7571);
  not g14071 (n_6750, n7572);
  and g14072 (n7573, n_6749, n_6750);
  not g14073 (n_6751, n7530);
  not g14074 (n_6752, n7573);
  and g14075 (n7574, n_6751, n_6752);
  and g14076 (n7575, n7530, n_6750);
  and g14077 (n7576, n_6749, n7575);
  not g14078 (n_6753, n7574);
  not g14079 (n_6754, n7576);
  and g14080 (n7577, n_6753, n_6754);
  not g14081 (n_6755, n7320);
  and g14082 (n7578, n_6755, n7577);
  not g14083 (n_6756, n7577);
  and g14084 (n7579, n7320, n_6756);
  not g14085 (n_6757, n7578);
  not g14086 (n_6758, n7579);
  and g14087 (n7580, n_6757, n_6758);
  and g14088 (n7581, n_6518, n_6521);
  not g14089 (n_6759, n7581);
  and g14090 (n7582, n_6517, n_6759);
  not g14091 (n_6760, n7580);
  and g14092 (n7583, n_6760, n7582);
  not g14093 (n_6761, n7582);
  and g14094 (n7584, n7580, n_6761);
  not g14095 (n_6762, n7583);
  not g14096 (n_6763, n7584);
  and g14097 (\asquared[57] , n_6762, n_6763);
  and g14098 (n7586, n_6748, n_6753);
  and g14099 (n7587, n_6742, n_6746);
  and g14100 (n7588, n_6651, n_6656);
  and g14101 (n7589, n_6618, n_6631);
  and g14102 (n7590, n7588, n7589);
  not g14103 (n_6764, n7588);
  not g14104 (n_6765, n7589);
  and g14105 (n7591, n_6764, n_6765);
  not g14106 (n_6766, n7590);
  not g14107 (n_6767, n7591);
  and g14108 (n7592, n_6766, n_6767);
  and g14109 (n7593, n_6586, n_6601);
  not g14110 (n_6768, n7592);
  and g14111 (n7594, n_6768, n7593);
  not g14112 (n_6769, n7593);
  and g14113 (n7595, n7592, n_6769);
  not g14114 (n_6770, n7594);
  not g14115 (n_6771, n7595);
  and g14116 (n7596, n_6770, n_6771);
  and g14117 (n7597, n_6604, n_6605);
  not g14118 (n_6772, n7597);
  and g14119 (n7598, n_6637, n_6772);
  not g14120 (n_6773, n7598);
  and g14121 (n7599, n7596, n_6773);
  not g14122 (n_6774, n7596);
  and g14123 (n7600, n_6774, n7598);
  not g14124 (n_6775, n7599);
  not g14125 (n_6776, n7600);
  and g14126 (n7601, n_6775, n_6776);
  and g14127 (n7602, n_6546, n_6561);
  and g14128 (n7603, n7359, n7390);
  not g14129 (n_6777, n7359);
  not g14130 (n_6778, n7390);
  and g14131 (n7604, n_6777, n_6778);
  not g14132 (n_6779, n7603);
  not g14133 (n_6780, n7604);
  and g14134 (n7605, n_6779, n_6780);
  not g14135 (n_6781, n7605);
  and g14136 (n7606, n7330, n_6781);
  not g14137 (n_6782, n7330);
  and g14138 (n7607, n_6782, n7605);
  not g14139 (n_6783, n7606);
  not g14140 (n_6784, n7607);
  and g14141 (n7608, n_6783, n_6784);
  and g14142 (n7609, n7375, n7444);
  not g14143 (n_6785, n7375);
  not g14144 (n_6786, n7444);
  and g14145 (n7610, n_6785, n_6786);
  not g14146 (n_6787, n7609);
  not g14147 (n_6788, n7610);
  and g14148 (n7611, n_6787, n_6788);
  and g14149 (n7612, n_6611, n_6614);
  not g14150 (n_6789, n7611);
  and g14151 (n7613, n_6789, n7612);
  not g14152 (n_6790, n7612);
  and g14153 (n7614, n7611, n_6790);
  not g14154 (n_6791, n7613);
  not g14155 (n_6792, n7614);
  and g14156 (n7615, n_6791, n_6792);
  and g14157 (n7616, n7608, n7615);
  not g14158 (n_6793, n7608);
  not g14159 (n_6794, n7615);
  and g14160 (n7617, n_6793, n_6794);
  not g14161 (n_6795, n7616);
  not g14162 (n_6796, n7617);
  and g14163 (n7618, n_6795, n_6796);
  not g14164 (n_6797, n7602);
  and g14165 (n7619, n_6797, n7618);
  not g14166 (n_6798, n7618);
  and g14167 (n7620, n7602, n_6798);
  not g14168 (n_6799, n7619);
  not g14169 (n_6800, n7620);
  and g14170 (n7621, n_6799, n_6800);
  and g14171 (n7622, n7601, n7621);
  not g14172 (n_6801, n7601);
  not g14173 (n_6802, n7621);
  and g14174 (n7623, n_6801, n_6802);
  not g14175 (n_6803, n7622);
  not g14176 (n_6804, n7623);
  and g14177 (n7624, n_6803, n_6804);
  not g14178 (n_6805, n7624);
  and g14179 (n7625, n7587, n_6805);
  not g14180 (n_6806, n7587);
  and g14181 (n7626, n_6806, n7624);
  not g14182 (n_6807, n7625);
  not g14183 (n_6808, n7626);
  and g14184 (n7627, n_6807, n_6808);
  and g14185 (n7628, n_6733, n_6738);
  and g14186 (n7629, n7409, n7543);
  not g14187 (n_6809, n7409);
  not g14188 (n_6810, n7543);
  and g14189 (n7630, n_6809, n_6810);
  not g14190 (n_6811, n7629);
  not g14191 (n_6812, n7630);
  and g14192 (n7631, n_6811, n_6812);
  not g14193 (n_6813, n7631);
  and g14194 (n7632, n7344, n_6813);
  not g14195 (n_6814, n7344);
  and g14196 (n7633, n_6814, n7631);
  not g14197 (n_6815, n7632);
  not g14198 (n_6816, n7633);
  and g14199 (n7634, n_6815, n_6816);
  and g14200 (n7635, n_6724, n_6730);
  not g14201 (n_6817, n7634);
  and g14202 (n7636, n_6817, n7635);
  not g14203 (n_6818, n7635);
  and g14204 (n7637, n7634, n_6818);
  not g14205 (n_6819, n7636);
  not g14206 (n_6820, n7637);
  and g14207 (n7638, n_6819, n_6820);
  and g14208 (n7639, \a[16] , \a[49] );
  and g14209 (n7640, n5620, n7639);
  and g14210 (n7641, n380, n6325);
  and g14211 (n7642, \a[16] , \a[50] );
  and g14212 (n7643, n5411, n7642);
  not g14213 (n_6821, n7641);
  not g14214 (n_6822, n7643);
  and g14215 (n7644, n_6821, n_6822);
  not g14216 (n_6823, n7640);
  not g14217 (n_6824, n7644);
  and g14218 (n7645, n_6823, n_6824);
  not g14219 (n_6825, n7645);
  and g14220 (n7646, n_6823, n_6825);
  and g14221 (n7647, \a[8] , \a[49] );
  and g14222 (n7648, \a[16] , \a[41] );
  not g14223 (n_6826, n7647);
  not g14224 (n_6827, n7648);
  and g14225 (n7649, n_6826, n_6827);
  not g14226 (n_6828, n7649);
  and g14227 (n7650, n7646, n_6828);
  and g14228 (n7651, \a[50] , n_6825);
  and g14229 (n7652, \a[7] , n7651);
  not g14230 (n_6829, n7650);
  not g14231 (n_6830, n7652);
  and g14232 (n7653, n_6829, n_6830);
  and g14233 (n7654, n1919, n3319);
  and g14234 (n7655, n1367, n4595);
  and g14235 (n7656, n1574, n3828);
  not g14236 (n_6831, n7655);
  not g14237 (n_6832, n7656);
  and g14238 (n7657, n_6831, n_6832);
  not g14239 (n_6833, n7654);
  not g14240 (n_6834, n7657);
  and g14241 (n7658, n_6833, n_6834);
  not g14242 (n_6835, n7658);
  and g14243 (n7659, \a[36] , n_6835);
  and g14244 (n7660, \a[21] , n7659);
  and g14245 (n7661, \a[22] , \a[35] );
  and g14246 (n7662, \a[23] , \a[34] );
  not g14247 (n_6836, n7661);
  not g14248 (n_6837, n7662);
  and g14249 (n7663, n_6836, n_6837);
  and g14250 (n7664, n_6833, n_6835);
  not g14251 (n_6838, n7663);
  and g14252 (n7665, n_6838, n7664);
  not g14253 (n_6839, n7660);
  not g14254 (n_6840, n7665);
  and g14255 (n7666, n_6839, n_6840);
  not g14256 (n_6841, n7653);
  not g14257 (n_6842, n7666);
  and g14258 (n7667, n_6841, n_6842);
  not g14259 (n_6843, n7667);
  and g14260 (n7668, n_6841, n_6843);
  and g14261 (n7669, n_6842, n_6843);
  not g14262 (n_6844, n7668);
  not g14263 (n_6845, n7669);
  and g14264 (n7670, n_6844, n_6845);
  and g14265 (n7671, n2463, n3812);
  and g14266 (n7672, n2301, n2598);
  and g14267 (n7673, n1904, n3143);
  not g14268 (n_6846, n7672);
  not g14269 (n_6847, n7673);
  and g14270 (n7674, n_6846, n_6847);
  not g14271 (n_6848, n7671);
  not g14272 (n_6849, n7674);
  and g14273 (n7675, n_6848, n_6849);
  not g14274 (n_6850, n7675);
  and g14275 (n7676, \a[33] , n_6850);
  and g14276 (n7677, \a[24] , n7676);
  and g14277 (n7678, n_6848, n_6850);
  and g14278 (n7679, \a[25] , \a[32] );
  and g14279 (n7680, \a[26] , \a[31] );
  not g14280 (n_6851, n7679);
  not g14281 (n_6852, n7680);
  and g14282 (n7681, n_6851, n_6852);
  not g14283 (n_6853, n7681);
  and g14284 (n7682, n7678, n_6853);
  not g14285 (n_6854, n7677);
  not g14286 (n_6855, n7682);
  and g14287 (n7683, n_6854, n_6855);
  not g14288 (n_6856, n7670);
  not g14289 (n_6857, n7683);
  and g14290 (n7684, n_6856, n_6857);
  not g14291 (n_6858, n7684);
  and g14292 (n7685, n_6856, n_6858);
  and g14293 (n7686, n_6857, n_6858);
  not g14294 (n_6859, n7685);
  not g14295 (n_6860, n7686);
  and g14296 (n7687, n_6859, n_6860);
  not g14297 (n_6861, n7687);
  and g14298 (n7688, n7638, n_6861);
  not g14299 (n_6862, n7638);
  and g14300 (n7689, n_6862, n7687);
  not g14301 (n_6863, n7628);
  not g14302 (n_6864, n7689);
  and g14303 (n7690, n_6863, n_6864);
  not g14304 (n_6865, n7688);
  and g14305 (n7691, n_6865, n7690);
  not g14306 (n_6866, n7691);
  and g14307 (n7692, n_6863, n_6866);
  and g14308 (n7693, n_6864, n_6866);
  and g14309 (n7694, n_6865, n7693);
  not g14310 (n_6867, n7692);
  not g14311 (n_6868, n7694);
  and g14312 (n7695, n_6867, n_6868);
  and g14313 (n7696, n_6693, n_6697);
  and g14314 (n7697, \a[53] , \a[55] );
  and g14315 (n7698, n252, n7697);
  and g14316 (n7699, \a[53] , \a[54] );
  and g14317 (n7700, n209, n7699);
  and g14318 (n7701, \a[54] , \a[55] );
  and g14319 (n7702, n218, n7701);
  not g14320 (n_6869, n7700);
  not g14321 (n_6870, n7702);
  and g14322 (n7703, n_6869, n_6870);
  not g14323 (n_6871, n7698);
  not g14324 (n_6872, n7703);
  and g14325 (n7704, n_6871, n_6872);
  not g14326 (n_6873, n7704);
  and g14327 (n7705, n_6871, n_6873);
  and g14328 (n7706, \a[2] , \a[55] );
  and g14329 (n7707, \a[4] , \a[53] );
  not g14330 (n_6874, n7706);
  not g14331 (n_6875, n7707);
  and g14332 (n7708, n_6874, n_6875);
  not g14333 (n_6876, n7708);
  and g14334 (n7709, n7705, n_6876);
  and g14335 (n7710, \a[54] , n_6873);
  and g14336 (n7711, \a[3] , n7710);
  not g14337 (n_6877, n7709);
  not g14338 (n_6878, n7711);
  and g14339 (n7712, n_6877, n_6878);
  and g14340 (n7713, \a[19] , \a[38] );
  and g14341 (n7714, \a[20] , \a[37] );
  not g14342 (n_6879, n7713);
  not g14343 (n_6880, n7714);
  and g14344 (n7715, n_6879, n_6880);
  and g14345 (n7716, n1490, n4565);
  not g14346 (n_6881, n7716);
  not g14349 (n_6882, n7715);
  not g14351 (n_6883, n7719);
  and g14352 (n7720, \a[52] , n_6883);
  and g14353 (n7721, \a[5] , n7720);
  and g14354 (n7722, n_6881, n_6883);
  and g14355 (n7723, n_6882, n7722);
  not g14356 (n_6884, n7721);
  not g14357 (n_6885, n7723);
  and g14358 (n7724, n_6884, n_6885);
  not g14359 (n_6886, n7712);
  not g14360 (n_6887, n7724);
  and g14361 (n7725, n_6886, n_6887);
  not g14362 (n_6888, n7725);
  and g14363 (n7726, n_6886, n_6888);
  and g14364 (n7727, n_6887, n_6888);
  not g14365 (n_6889, n7726);
  not g14366 (n_6890, n7727);
  and g14367 (n7728, n_6889, n_6890);
  and g14368 (n7729, \a[9] , \a[48] );
  and g14369 (n7730, \a[10] , \a[47] );
  not g14370 (n_6891, n7729);
  not g14371 (n_6892, n7730);
  and g14372 (n7731, n_6891, n_6892);
  and g14373 (n7732, n484, n6252);
  not g14374 (n_6893, n7732);
  not g14377 (n_6894, n7731);
  not g14379 (n_6895, n7735);
  and g14380 (n7736, \a[42] , n_6895);
  and g14381 (n7737, \a[15] , n7736);
  and g14382 (n7738, n_6893, n_6895);
  and g14383 (n7739, n_6894, n7738);
  not g14384 (n_6896, n7737);
  not g14385 (n_6897, n7739);
  and g14386 (n7740, n_6896, n_6897);
  not g14387 (n_6898, n7728);
  not g14388 (n_6899, n7740);
  and g14389 (n7741, n_6898, n_6899);
  not g14390 (n_6900, n7741);
  and g14391 (n7742, n_6898, n_6900);
  and g14392 (n7743, n_6899, n_6900);
  not g14393 (n_6901, n7742);
  not g14394 (n_6902, n7743);
  and g14395 (n7744, n_6901, n_6902);
  and g14396 (n7745, \a[11] , \a[46] );
  not g14397 (n_6903, n6168);
  not g14398 (n_6904, n7745);
  and g14399 (n7746, n_6903, n_6904);
  and g14400 (n7747, \a[44] , \a[46] );
  and g14401 (n7748, n818, n7747);
  and g14402 (n7749, n745, n5296);
  and g14403 (n7750, n6933, n7400);
  not g14404 (n_6905, n7749);
  not g14405 (n_6906, n7750);
  and g14406 (n7751, n_6905, n_6906);
  not g14407 (n_6907, n7748);
  not g14408 (n_6908, n7751);
  and g14409 (n7752, n_6907, n_6908);
  not g14410 (n_6909, n7752);
  and g14411 (n7753, n_6907, n_6909);
  not g14412 (n_6910, n7746);
  and g14413 (n7754, n_6910, n7753);
  and g14414 (n7755, \a[43] , n_6909);
  and g14415 (n7756, \a[14] , n7755);
  not g14416 (n_6911, n7754);
  not g14417 (n_6912, n7756);
  and g14418 (n7757, n_6911, n_6912);
  not g14419 (n_6913, n2334);
  not g14420 (n_6914, n2922);
  and g14421 (n7758, n_6913, n_6914);
  and g14422 (n7759, n2331, n2617);
  not g14423 (n_6915, n7759);
  not g14426 (n_6916, n7758);
  not g14428 (n_6917, n7762);
  and g14429 (n7763, \a[45] , n_6917);
  and g14430 (n7764, \a[12] , n7763);
  and g14431 (n7765, n_6915, n_6917);
  and g14432 (n7766, n_6916, n7765);
  not g14433 (n_6918, n7764);
  not g14434 (n_6919, n7766);
  and g14435 (n7767, n_6918, n_6919);
  not g14436 (n_6920, n7757);
  not g14437 (n_6921, n7767);
  and g14438 (n7768, n_6920, n_6921);
  not g14439 (n_6922, n7768);
  and g14440 (n7769, n_6920, n_6922);
  and g14441 (n7770, n_6921, n_6922);
  not g14442 (n_6923, n7769);
  not g14443 (n_6924, n7770);
  and g14444 (n7771, n_6923, n_6924);
  and g14445 (n7772, \a[17] , \a[51] );
  and g14446 (n7773, n4972, n7772);
  and g14447 (n7774, \a[39] , \a[51] );
  and g14448 (n7775, n1478, n7774);
  and g14449 (n7776, n1052, n4171);
  not g14450 (n_6925, n7775);
  not g14451 (n_6926, n7776);
  and g14452 (n7777, n_6925, n_6926);
  not g14453 (n_6927, n7773);
  not g14454 (n_6928, n7777);
  and g14455 (n7778, n_6927, n_6928);
  not g14456 (n_6929, n7778);
  and g14457 (n7779, \a[39] , n_6929);
  and g14458 (n7780, \a[18] , n7779);
  and g14459 (n7781, n_6927, n_6929);
  and g14460 (n7782, \a[6] , \a[51] );
  and g14461 (n7783, \a[17] , \a[40] );
  not g14462 (n_6930, n7782);
  not g14463 (n_6931, n7783);
  and g14464 (n7784, n_6930, n_6931);
  not g14465 (n_6932, n7784);
  and g14466 (n7785, n7781, n_6932);
  not g14467 (n_6933, n7780);
  not g14468 (n_6934, n7785);
  and g14469 (n7786, n_6933, n_6934);
  not g14470 (n_6935, n7771);
  not g14471 (n_6936, n7786);
  and g14472 (n7787, n_6935, n_6936);
  not g14473 (n_6937, n7787);
  and g14474 (n7788, n_6935, n_6937);
  and g14475 (n7789, n_6936, n_6937);
  not g14476 (n_6938, n7788);
  not g14477 (n_6939, n7789);
  and g14478 (n7790, n_6938, n_6939);
  and g14479 (n7791, n7744, n7790);
  not g14480 (n_6940, n7744);
  not g14481 (n_6941, n7790);
  and g14482 (n7792, n_6940, n_6941);
  not g14483 (n_6942, n7791);
  not g14484 (n_6943, n7792);
  and g14485 (n7793, n_6942, n_6943);
  not g14486 (n_6944, n7696);
  and g14487 (n7794, n_6944, n7793);
  not g14488 (n_6945, n7793);
  and g14489 (n7795, n7696, n_6945);
  not g14490 (n_6946, n7794);
  not g14491 (n_6947, n7795);
  and g14492 (n7796, n_6946, n_6947);
  and g14493 (n7797, n7695, n7796);
  not g14494 (n_6948, n7695);
  not g14495 (n_6949, n7796);
  and g14496 (n7798, n_6948, n_6949);
  not g14497 (n_6950, n7797);
  not g14498 (n_6951, n7798);
  and g14499 (n7799, n_6950, n_6951);
  not g14500 (n_6952, n7799);
  and g14501 (n7800, n7627, n_6952);
  not g14502 (n_6953, n7800);
  and g14503 (n7801, n7627, n_6953);
  and g14504 (n7802, n_6952, n_6953);
  not g14505 (n_6954, n7801);
  not g14506 (n_6955, n7802);
  and g14507 (n7803, n_6954, n_6955);
  and g14508 (n7804, n_6707, n_6712);
  and g14509 (n7805, n_6667, n_6671);
  and g14510 (n7806, n_6699, n_6704);
  and g14511 (n7807, n_6685, n_6689);
  and g14512 (n7808, n_6660, n_6664);
  and g14513 (n7809, n7807, n7808);
  not g14514 (n_6956, n7807);
  not g14515 (n_6957, n7808);
  and g14516 (n7810, n_6956, n_6957);
  not g14517 (n_6958, n7809);
  not g14518 (n_6959, n7810);
  and g14519 (n7811, n_6958, n_6959);
  and g14520 (n7812, \a[0] , \a[57] );
  and g14521 (n7813, n7465, n7812);
  not g14522 (n_6961, n7813);
  and g14523 (n7814, n7465, n_6961);
  and g14524 (n7815, n_6649, n7812);
  not g14525 (n_6962, n7814);
  not g14526 (n_6963, n7815);
  and g14527 (n7816, n_6962, n_6963);
  and g14528 (n7817, \a[1] , \a[56] );
  and g14529 (n7818, \a[29] , n7817);
  not g14530 (n_6964, n7818);
  and g14531 (n7819, \a[29] , n_6964);
  and g14532 (n7820, n7817, n_6964);
  not g14533 (n_6965, n7819);
  not g14534 (n_6966, n7820);
  and g14535 (n7821, n_6965, n_6966);
  not g14536 (n_6967, n7816);
  not g14537 (n_6968, n7821);
  and g14538 (n7822, n_6967, n_6968);
  not g14539 (n_6969, n7822);
  and g14540 (n7823, n_6967, n_6969);
  and g14541 (n7824, n_6968, n_6969);
  not g14542 (n_6970, n7823);
  not g14543 (n_6971, n7824);
  and g14544 (n7825, n_6970, n_6971);
  and g14545 (n7826, n_6641, n_6645);
  and g14546 (n7827, n7825, n7826);
  not g14547 (n_6972, n7825);
  not g14548 (n_6973, n7826);
  and g14549 (n7828, n_6972, n_6973);
  not g14550 (n_6974, n7827);
  not g14551 (n_6975, n7828);
  and g14552 (n7829, n_6974, n_6975);
  and g14553 (n7830, n_6677, n_6681);
  not g14554 (n_6976, n7829);
  and g14555 (n7831, n_6976, n7830);
  not g14556 (n_6977, n7830);
  and g14557 (n7832, n7829, n_6977);
  not g14558 (n_6978, n7831);
  not g14559 (n_6979, n7832);
  and g14560 (n7833, n_6978, n_6979);
  and g14561 (n7834, n7811, n7833);
  not g14562 (n_6980, n7811);
  not g14563 (n_6981, n7833);
  and g14564 (n7835, n_6980, n_6981);
  not g14565 (n_6982, n7834);
  not g14566 (n_6983, n7835);
  and g14567 (n7836, n_6982, n_6983);
  not g14568 (n_6984, n7806);
  and g14569 (n7837, n_6984, n7836);
  not g14570 (n_6985, n7836);
  and g14571 (n7838, n7806, n_6985);
  not g14572 (n_6986, n7837);
  not g14573 (n_6987, n7838);
  and g14574 (n7839, n_6986, n_6987);
  not g14575 (n_6988, n7805);
  and g14576 (n7840, n_6988, n7839);
  not g14577 (n_6989, n7839);
  and g14578 (n7841, n7805, n_6989);
  not g14579 (n_6990, n7840);
  not g14580 (n_6991, n7841);
  and g14581 (n7842, n_6990, n_6991);
  not g14582 (n_6992, n7804);
  and g14583 (n7843, n_6992, n7842);
  not g14584 (n_6993, n7843);
  and g14585 (n7844, n_6992, n_6993);
  and g14586 (n7845, n7842, n_6993);
  not g14587 (n_6994, n7844);
  not g14588 (n_6995, n7845);
  and g14589 (n7846, n_6994, n_6995);
  not g14590 (n_6996, n7803);
  not g14591 (n_6997, n7846);
  and g14592 (n7847, n_6996, n_6997);
  and g14593 (n7848, n7803, n_6995);
  and g14594 (n7849, n_6994, n7848);
  not g14595 (n_6998, n7847);
  not g14596 (n_6999, n7849);
  and g14597 (n7850, n_6998, n_6999);
  not g14598 (n_7000, n7586);
  and g14599 (n7851, n_7000, n7850);
  not g14600 (n_7001, n7850);
  and g14601 (n7852, n7586, n_7001);
  not g14602 (n_7002, n7851);
  not g14603 (n_7003, n7852);
  and g14604 (n7853, n_7002, n_7003);
  and g14605 (n7854, n_6758, n_6761);
  not g14606 (n_7004, n7854);
  and g14607 (n7855, n_6757, n_7004);
  not g14608 (n_7005, n7853);
  and g14609 (n7856, n_7005, n7855);
  not g14610 (n_7006, n7855);
  and g14611 (n7857, n7853, n_7006);
  not g14612 (n_7007, n7856);
  not g14613 (n_7008, n7857);
  and g14614 (\asquared[58] , n_7007, n_7008);
  and g14615 (n7859, n_7003, n_7006);
  not g14616 (n_7009, n7859);
  and g14617 (n7860, n_7002, n_7009);
  and g14618 (n7861, n_6993, n_6998);
  and g14619 (n7862, n_6808, n_6953);
  and g14620 (n7863, n_6775, n_6803);
  and g14621 (n7864, n_6820, n_6865);
  and g14622 (n7865, n_6812, n_6816);
  and g14623 (n7866, n_6788, n_6792);
  and g14624 (n7867, n7865, n7866);
  not g14625 (n_7010, n7865);
  not g14626 (n_7011, n7866);
  and g14627 (n7868, n_7010, n_7011);
  not g14628 (n_7012, n7867);
  not g14629 (n_7013, n7868);
  and g14630 (n7869, n_7012, n_7013);
  and g14631 (n7870, n_6780, n_6784);
  not g14632 (n_7014, n7869);
  and g14633 (n7871, n_7014, n7870);
  not g14634 (n_7015, n7870);
  and g14635 (n7872, n7869, n_7015);
  not g14636 (n_7016, n7871);
  not g14637 (n_7017, n7872);
  and g14638 (n7873, n_7016, n_7017);
  and g14639 (n7874, n_6795, n_6799);
  not g14640 (n_7018, n7874);
  and g14641 (n7875, n7873, n_7018);
  not g14642 (n_7019, n7873);
  and g14643 (n7876, n_7019, n7874);
  not g14644 (n_7020, n7875);
  not g14645 (n_7021, n7876);
  and g14646 (n7877, n_7020, n_7021);
  not g14647 (n_7022, n7864);
  and g14648 (n7878, n_7022, n7877);
  not g14649 (n_7023, n7877);
  and g14650 (n7879, n7864, n_7023);
  not g14651 (n_7024, n7878);
  not g14652 (n_7025, n7879);
  and g14653 (n7880, n_7024, n_7025);
  not g14654 (n_7026, n7880);
  and g14655 (n7881, n7863, n_7026);
  not g14656 (n_7027, n7863);
  and g14657 (n7882, n_7027, n7880);
  not g14658 (n_7028, n7881);
  not g14659 (n_7029, n7882);
  and g14660 (n7883, n_7028, n_7029);
  and g14661 (n7884, n_6948, n7796);
  not g14662 (n_7030, n7884);
  and g14663 (n7885, n_6866, n_7030);
  not g14664 (n_7031, n7885);
  and g14665 (n7886, n7883, n_7031);
  not g14666 (n_7032, n7883);
  and g14667 (n7887, n_7032, n7885);
  not g14668 (n_7033, n7886);
  not g14669 (n_7034, n7887);
  and g14670 (n7888, n_7033, n_7034);
  not g14671 (n_7035, n7888);
  and g14672 (n7889, n7862, n_7035);
  not g14673 (n_7036, n7862);
  and g14674 (n7890, n_7036, n7888);
  not g14675 (n_7037, n7889);
  not g14676 (n_7038, n7890);
  and g14677 (n7891, n_7037, n_7038);
  and g14678 (n7892, n_6986, n_6990);
  and g14679 (n7893, n_6943, n_6946);
  and g14680 (n7894, n_6922, n_6937);
  and g14681 (n7895, n_6888, n_6900);
  and g14682 (n7896, \a[1] , \a[57] );
  and g14683 (n7897, n3110, n7896);
  not g14684 (n_7039, n3110);
  not g14685 (n_7040, n7896);
  and g14686 (n7898, n_7039, n_7040);
  not g14687 (n_7041, n7897);
  not g14688 (n_7042, n7898);
  and g14689 (n7899, n_7041, n_7042);
  not g14690 (n_7043, n7899);
  and g14691 (n7900, n_6964, n_7043);
  and g14692 (n7901, n7818, n7899);
  not g14693 (n_7044, n7900);
  not g14694 (n_7045, n7901);
  and g14695 (n7902, n_7044, n_7045);
  not g14696 (n_7046, n7765);
  and g14697 (n7903, n_7046, n7902);
  not g14698 (n_7047, n7902);
  and g14699 (n7904, n7765, n_7047);
  not g14700 (n_7048, n7903);
  not g14701 (n_7049, n7904);
  and g14702 (n7905, n_7048, n_7049);
  not g14703 (n_7050, n7895);
  and g14704 (n7906, n_7050, n7905);
  not g14705 (n_7051, n7906);
  and g14706 (n7907, n_7050, n_7051);
  and g14707 (n7908, n7905, n_7051);
  not g14708 (n_7052, n7907);
  not g14709 (n_7053, n7908);
  and g14710 (n7909, n_7052, n_7053);
  not g14711 (n_7054, n7894);
  not g14712 (n_7055, n7909);
  and g14713 (n7910, n_7054, n_7055);
  and g14714 (n7911, n7894, n_7053);
  and g14715 (n7912, n_7052, n7911);
  not g14716 (n_7056, n7910);
  not g14717 (n_7057, n7912);
  and g14718 (n7913, n_7056, n_7057);
  not g14719 (n_7058, n7893);
  and g14720 (n7914, n_7058, n7913);
  not g14721 (n_7059, n7913);
  and g14722 (n7915, n7893, n_7059);
  not g14723 (n_7060, n7914);
  not g14724 (n_7061, n7915);
  and g14725 (n7916, n_7060, n_7061);
  and g14726 (n7917, n_6843, n_6858);
  and g14727 (n7918, n7678, n7738);
  not g14728 (n_7062, n7678);
  not g14729 (n_7063, n7738);
  and g14730 (n7919, n_7062, n_7063);
  not g14731 (n_7064, n7918);
  not g14732 (n_7065, n7919);
  and g14733 (n7920, n_7064, n_7065);
  not g14734 (n_7066, n7920);
  and g14735 (n7921, n7664, n_7066);
  not g14736 (n_7067, n7664);
  and g14737 (n7922, n_7067, n7920);
  not g14738 (n_7068, n7921);
  not g14739 (n_7069, n7922);
  and g14740 (n7923, n_7068, n_7069);
  and g14741 (n7924, n7705, n7722);
  not g14742 (n_7070, n7705);
  not g14743 (n_7071, n7722);
  and g14744 (n7925, n_7070, n_7071);
  not g14745 (n_7072, n7924);
  not g14746 (n_7073, n7925);
  and g14747 (n7926, n_7072, n_7073);
  not g14748 (n_7074, n7926);
  and g14749 (n7927, n7753, n_7074);
  not g14750 (n_7075, n7753);
  and g14751 (n7928, n_7075, n7926);
  not g14752 (n_7076, n7927);
  not g14753 (n_7077, n7928);
  and g14754 (n7929, n_7076, n_7077);
  and g14755 (n7930, n7923, n7929);
  not g14756 (n_7078, n7923);
  not g14757 (n_7079, n7929);
  and g14758 (n7931, n_7078, n_7079);
  not g14759 (n_7080, n7930);
  not g14760 (n_7081, n7931);
  and g14761 (n7932, n_7080, n_7081);
  not g14762 (n_7082, n7917);
  and g14763 (n7933, n_7082, n7932);
  not g14764 (n_7083, n7932);
  and g14765 (n7934, n7917, n_7083);
  not g14766 (n_7084, n7933);
  not g14767 (n_7085, n7934);
  and g14768 (n7935, n_7084, n_7085);
  and g14769 (n7936, n7916, n7935);
  not g14770 (n_7086, n7916);
  not g14771 (n_7087, n7935);
  and g14772 (n7937, n_7086, n_7087);
  not g14773 (n_7088, n7936);
  not g14774 (n_7089, n7937);
  and g14775 (n7938, n_7088, n_7089);
  not g14776 (n_7090, n7938);
  and g14777 (n7939, n7892, n_7090);
  not g14778 (n_7091, n7892);
  and g14779 (n7940, n_7091, n7938);
  not g14780 (n_7092, n7939);
  not g14781 (n_7093, n7940);
  and g14782 (n7941, n_7092, n_7093);
  and g14783 (n7942, \a[56] , \a[58] );
  and g14784 (n7943, n196, n7942);
  and g14785 (n7944, n252, n7421);
  not g14786 (n_7095, n7943);
  not g14787 (n_7096, n7944);
  and g14788 (n7945, n_7095, n_7096);
  and g14789 (n7946, \a[0] , \a[58] );
  and g14790 (n7947, \a[4] , \a[54] );
  and g14791 (n7948, n7946, n7947);
  not g14792 (n_7097, n7945);
  not g14793 (n_7098, n7948);
  and g14794 (n7949, n_7097, n_7098);
  not g14795 (n_7099, n7949);
  and g14796 (n7950, n_7098, n_7099);
  not g14797 (n_7100, n7946);
  not g14798 (n_7101, n7947);
  and g14799 (n7951, n_7100, n_7101);
  not g14800 (n_7102, n7951);
  and g14801 (n7952, n7950, n_7102);
  and g14802 (n7953, \a[2] , \a[56] );
  and g14803 (n7954, n_7099, n7953);
  not g14804 (n_7103, n7952);
  not g14805 (n_7104, n7954);
  and g14806 (n7955, n_7103, n_7104);
  and g14807 (n7956, \a[20] , \a[38] );
  and g14808 (n7957, \a[21] , \a[37] );
  not g14809 (n_7105, n7956);
  not g14810 (n_7106, n7957);
  and g14811 (n7958, n_7105, n_7106);
  and g14812 (n7959, n1494, n4565);
  not g14813 (n_7107, n7959);
  not g14816 (n_7108, n7958);
  not g14818 (n_7109, n7962);
  and g14819 (n7963, \a[53] , n_7109);
  and g14820 (n7964, \a[5] , n7963);
  and g14821 (n7965, n_7107, n_7109);
  and g14822 (n7966, n_7108, n7965);
  not g14823 (n_7110, n7964);
  not g14824 (n_7111, n7966);
  and g14825 (n7967, n_7110, n_7111);
  not g14826 (n_7112, n7955);
  not g14827 (n_7113, n7967);
  and g14828 (n7968, n_7112, n_7113);
  not g14829 (n_7114, n7968);
  and g14830 (n7969, n_7112, n_7114);
  and g14831 (n7970, n_7113, n_7114);
  not g14832 (n_7115, n7969);
  not g14833 (n_7116, n7970);
  and g14834 (n7971, n_7115, n_7116);
  and g14835 (n7972, \a[42] , \a[49] );
  and g14836 (n7973, n847, n7972);
  and g14837 (n7974, n1048, n5344);
  and g14838 (n7975, n5956, n7063);
  not g14839 (n_7117, n7974);
  not g14840 (n_7118, n7975);
  and g14841 (n7976, n_7117, n_7118);
  not g14842 (n_7119, n7973);
  not g14843 (n_7120, n7976);
  and g14844 (n7977, n_7119, n_7120);
  not g14845 (n_7121, n7977);
  and g14846 (n7978, \a[41] , n_7121);
  and g14847 (n7979, \a[17] , n7978);
  and g14848 (n7980, \a[9] , \a[49] );
  and g14849 (n7981, \a[16] , \a[42] );
  not g14850 (n_7122, n7980);
  not g14851 (n_7123, n7981);
  and g14852 (n7982, n_7122, n_7123);
  and g14853 (n7983, n_7119, n_7121);
  not g14854 (n_7124, n7982);
  and g14855 (n7984, n_7124, n7983);
  not g14856 (n_7125, n7979);
  not g14857 (n_7126, n7984);
  and g14858 (n7985, n_7125, n_7126);
  not g14859 (n_7127, n7971);
  not g14860 (n_7128, n7985);
  and g14861 (n7986, n_7127, n_7128);
  not g14862 (n_7129, n7986);
  and g14863 (n7987, n_7127, n_7129);
  and g14864 (n7988, n_7128, n_7129);
  not g14865 (n_7130, n7987);
  not g14866 (n_7131, n7988);
  and g14867 (n7989, n_7130, n_7131);
  and g14868 (n7990, \a[7] , \a[51] );
  and g14869 (n7991, \a[8] , \a[50] );
  not g14870 (n_7132, n7990);
  not g14871 (n_7133, n7991);
  and g14872 (n7992, n_7132, n_7133);
  and g14873 (n7993, n380, n6564);
  not g14874 (n_7134, n7993);
  not g14877 (n_7135, n7992);
  not g14879 (n_7136, n7996);
  and g14880 (n7997, n_7134, n_7136);
  and g14881 (n7998, n_7135, n7997);
  and g14882 (n7999, \a[40] , n_7136);
  and g14883 (n8000, \a[18] , n7999);
  not g14884 (n_7137, n7998);
  not g14885 (n_7138, n8000);
  and g14886 (n8001, n_7137, n_7138);
  and g14887 (n8002, n1666, n3319);
  and g14888 (n8003, n2115, n4595);
  and g14889 (n8004, n1919, n3828);
  not g14890 (n_7139, n8003);
  not g14891 (n_7140, n8004);
  and g14892 (n8005, n_7139, n_7140);
  not g14893 (n_7141, n8002);
  not g14894 (n_7142, n8005);
  and g14895 (n8006, n_7141, n_7142);
  not g14896 (n_7143, n8006);
  and g14897 (n8007, \a[36] , n_7143);
  and g14898 (n8008, \a[22] , n8007);
  and g14899 (n8009, n_7141, n_7143);
  and g14900 (n8010, \a[23] , \a[35] );
  and g14901 (n8011, \a[24] , \a[34] );
  not g14902 (n_7144, n8010);
  not g14903 (n_7145, n8011);
  and g14904 (n8012, n_7144, n_7145);
  not g14905 (n_7146, n8012);
  and g14906 (n8013, n8009, n_7146);
  not g14907 (n_7147, n8008);
  not g14908 (n_7148, n8013);
  and g14909 (n8014, n_7147, n_7148);
  not g14910 (n_7149, n8001);
  not g14911 (n_7150, n8014);
  and g14912 (n8015, n_7149, n_7150);
  not g14913 (n_7151, n8015);
  and g14914 (n8016, n_7149, n_7151);
  and g14915 (n8017, n_7150, n_7151);
  not g14916 (n_7152, n8016);
  not g14917 (n_7153, n8017);
  and g14918 (n8018, n_7152, n_7153);
  and g14919 (n8019, n2227, n3812);
  and g14920 (n8020, n2598, n2633);
  and g14921 (n8021, n2463, n3143);
  not g14922 (n_7154, n8020);
  not g14923 (n_7155, n8021);
  and g14924 (n8022, n_7154, n_7155);
  not g14925 (n_7156, n8019);
  not g14926 (n_7157, n8022);
  and g14927 (n8023, n_7156, n_7157);
  not g14928 (n_7158, n8023);
  and g14929 (n8024, n3301, n_7158);
  and g14930 (n8025, n_7156, n_7158);
  and g14931 (n8026, \a[27] , \a[31] );
  not g14932 (n_7159, n3266);
  not g14933 (n_7160, n8026);
  and g14934 (n8027, n_7159, n_7160);
  not g14935 (n_7161, n8027);
  and g14936 (n8028, n8025, n_7161);
  not g14937 (n_7162, n8024);
  not g14938 (n_7163, n8028);
  and g14939 (n8029, n_7162, n_7163);
  not g14940 (n_7164, n8018);
  not g14941 (n_7165, n8029);
  and g14942 (n8030, n_7164, n_7165);
  not g14943 (n_7166, n8030);
  and g14944 (n8031, n_7164, n_7166);
  and g14945 (n8032, n_7165, n_7166);
  not g14946 (n_7167, n8031);
  not g14947 (n_7168, n8032);
  and g14948 (n8033, n_7167, n_7168);
  not g14949 (n_7169, n7989);
  and g14950 (n8034, n_7169, n8033);
  not g14951 (n_7170, n8033);
  and g14952 (n8035, n7989, n_7170);
  not g14953 (n_7171, n8034);
  not g14954 (n_7172, n8035);
  and g14955 (n8036, n_7171, n_7172);
  and g14956 (n8037, n_6767, n_6771);
  and g14957 (n8038, n8036, n8037);
  not g14958 (n_7173, n8036);
  not g14959 (n_7174, n8037);
  and g14960 (n8039, n_7173, n_7174);
  not g14961 (n_7175, n8038);
  not g14962 (n_7176, n8039);
  and g14963 (n8040, n_7175, n_7176);
  and g14964 (n8041, n_6959, n_6982);
  and g14965 (n8042, n7646, n7781);
  not g14966 (n_7177, n7646);
  not g14967 (n_7178, n7781);
  and g14968 (n8043, n_7177, n_7178);
  not g14969 (n_7179, n8042);
  not g14970 (n_7180, n8043);
  and g14971 (n8044, n_7179, n_7180);
  and g14972 (n8045, n_6961, n_6969);
  not g14973 (n_7181, n8044);
  and g14974 (n8046, n_7181, n8045);
  not g14975 (n_7182, n8045);
  and g14976 (n8047, n8044, n_7182);
  not g14977 (n_7183, n8046);
  not g14978 (n_7184, n8047);
  and g14979 (n8048, n_7183, n_7184);
  and g14980 (n8049, n_6975, n_6979);
  not g14981 (n_7185, n8048);
  and g14982 (n8050, n_7185, n8049);
  not g14983 (n_7186, n8049);
  and g14984 (n8051, n8048, n_7186);
  not g14985 (n_7187, n8050);
  not g14986 (n_7188, n8051);
  and g14987 (n8052, n_7187, n_7188);
  and g14988 (n8053, \a[43] , \a[47] );
  and g14989 (n8054, n816, n8053);
  and g14990 (n8055, n723, n6252);
  and g14991 (n8056, n6659, n7351);
  not g14992 (n_7189, n8055);
  not g14993 (n_7190, n8056);
  and g14994 (n8057, n_7189, n_7190);
  not g14995 (n_7191, n8054);
  not g14996 (n_7192, n8057);
  and g14997 (n8058, n_7191, n_7192);
  not g14998 (n_7193, n8058);
  and g14999 (n8059, n_7191, n_7193);
  and g15000 (n8060, \a[11] , \a[47] );
  not g15001 (n_7194, n5647);
  not g15002 (n_7195, n8060);
  and g15003 (n8061, n_7194, n_7195);
  not g15004 (n_7196, n8061);
  and g15005 (n8062, n8059, n_7196);
  and g15006 (n8063, \a[48] , n_7193);
  and g15007 (n8064, \a[10] , n8063);
  not g15008 (n_7197, n8062);
  not g15009 (n_7198, n8064);
  and g15010 (n8065, n_7197, n_7198);
  and g15011 (n8066, n748, n5560);
  and g15012 (n8067, n606, n7747);
  and g15013 (n8068, n745, n5713);
  not g15014 (n_7199, n8067);
  not g15015 (n_7200, n8068);
  and g15016 (n8069, n_7199, n_7200);
  not g15017 (n_7201, n8066);
  not g15018 (n_7202, n8069);
  and g15019 (n8070, n_7201, n_7202);
  not g15020 (n_7203, n8070);
  and g15021 (n8071, n6621, n_7203);
  and g15022 (n8072, n_7201, n_7203);
  and g15023 (n8073, \a[12] , \a[46] );
  not g15024 (n_7204, n7186);
  not g15025 (n_7205, n8073);
  and g15026 (n8074, n_7204, n_7205);
  not g15027 (n_7206, n8074);
  and g15028 (n8075, n8072, n_7206);
  not g15029 (n_7207, n8071);
  not g15030 (n_7208, n8075);
  and g15031 (n8076, n_7207, n_7208);
  not g15032 (n_7209, n8065);
  not g15033 (n_7210, n8076);
  and g15034 (n8077, n_7209, n_7210);
  not g15035 (n_7211, n8077);
  and g15036 (n8078, n_7209, n_7211);
  and g15037 (n8079, n_7210, n_7211);
  not g15038 (n_7212, n8078);
  not g15039 (n_7213, n8079);
  and g15040 (n8080, n_7212, n_7213);
  and g15041 (n8081, \a[6] , \a[52] );
  and g15042 (n8082, \a[19] , \a[39] );
  not g15043 (n_7214, n8081);
  not g15044 (n_7215, n8082);
  and g15045 (n8083, n_7214, n_7215);
  and g15046 (n8084, n8081, n8082);
  not g15047 (n_7216, n8084);
  not g15050 (n_7217, n8083);
  not g15052 (n_7218, n8087);
  and g15053 (n8088, \a[55] , n_7218);
  and g15054 (n8089, \a[3] , n8088);
  and g15055 (n8090, n_7216, n_7218);
  and g15056 (n8091, n_7217, n8090);
  not g15057 (n_7219, n8089);
  not g15058 (n_7220, n8091);
  and g15059 (n8092, n_7219, n_7220);
  not g15060 (n_7221, n8080);
  not g15061 (n_7222, n8092);
  and g15062 (n8093, n_7221, n_7222);
  not g15063 (n_7223, n8093);
  and g15064 (n8094, n_7221, n_7223);
  and g15065 (n8095, n_7222, n_7223);
  not g15066 (n_7224, n8094);
  not g15067 (n_7225, n8095);
  and g15068 (n8096, n_7224, n_7225);
  not g15069 (n_7226, n8052);
  and g15070 (n8097, n_7226, n8096);
  not g15071 (n_7227, n8096);
  and g15072 (n8098, n8052, n_7227);
  not g15073 (n_7228, n8097);
  not g15074 (n_7229, n8098);
  and g15075 (n8099, n_7228, n_7229);
  not g15076 (n_7230, n8041);
  and g15077 (n8100, n_7230, n8099);
  not g15078 (n_7231, n8100);
  and g15079 (n8101, n_7230, n_7231);
  and g15080 (n8102, n8099, n_7231);
  not g15081 (n_7232, n8101);
  not g15082 (n_7233, n8102);
  and g15083 (n8103, n_7232, n_7233);
  not g15084 (n_7234, n8103);
  and g15085 (n8104, n8040, n_7234);
  not g15086 (n_7235, n8104);
  and g15087 (n8105, n8040, n_7235);
  and g15088 (n8106, n_7234, n_7235);
  not g15089 (n_7236, n8105);
  not g15090 (n_7237, n8106);
  and g15091 (n8107, n_7236, n_7237);
  not g15092 (n_7238, n8107);
  and g15093 (n8108, n7941, n_7238);
  not g15094 (n_7239, n8108);
  and g15095 (n8109, n7941, n_7239);
  and g15096 (n8110, n_7238, n_7239);
  not g15097 (n_7240, n8109);
  not g15098 (n_7241, n8110);
  and g15099 (n8111, n_7240, n_7241);
  not g15100 (n_7242, n7891);
  and g15101 (n8112, n_7242, n8111);
  not g15102 (n_7243, n8111);
  and g15103 (n8113, n7891, n_7243);
  not g15104 (n_7244, n8112);
  not g15105 (n_7245, n8113);
  and g15106 (n8114, n_7244, n_7245);
  not g15107 (n_7246, n7861);
  and g15108 (n8115, n_7246, n8114);
  not g15109 (n_7247, n8114);
  and g15110 (n8116, n7861, n_7247);
  not g15111 (n_7248, n8115);
  not g15112 (n_7249, n8116);
  and g15113 (n8117, n_7248, n_7249);
  not g15114 (n_7250, n8117);
  and g15115 (n8118, n7860, n_7250);
  not g15116 (n_7251, n7860);
  and g15117 (n8119, n_7251, n_7249);
  and g15118 (n8120, n_7248, n8119);
  not g15119 (n_7252, n8118);
  not g15120 (n_7253, n8120);
  and g15121 (\asquared[59] , n_7252, n_7253);
  and g15122 (n8122, n_7093, n_7239);
  and g15123 (n8123, n_7231, n_7235);
  and g15124 (n8124, n_7060, n_7088);
  and g15125 (n8125, n_7188, n_7229);
  and g15126 (n8126, n_7180, n_7184);
  and g15127 (n8127, n_7073, n_7077);
  and g15128 (n8128, n8126, n8127);
  not g15129 (n_7254, n8126);
  not g15130 (n_7255, n8127);
  and g15131 (n8129, n_7254, n_7255);
  not g15132 (n_7256, n8128);
  not g15133 (n_7257, n8129);
  and g15134 (n8130, n_7256, n_7257);
  and g15135 (n8131, n_7065, n_7069);
  not g15136 (n_7258, n8130);
  and g15137 (n8132, n_7258, n8131);
  not g15138 (n_7259, n8131);
  and g15139 (n8133, n8130, n_7259);
  not g15140 (n_7260, n8132);
  not g15141 (n_7261, n8133);
  and g15142 (n8134, n_7260, n_7261);
  and g15143 (n8135, n_7080, n_7084);
  not g15144 (n_7262, n8135);
  and g15145 (n8136, n8134, n_7262);
  not g15146 (n_7263, n8134);
  and g15147 (n8137, n_7263, n8135);
  not g15148 (n_7264, n8136);
  not g15149 (n_7265, n8137);
  and g15150 (n8138, n_7264, n_7265);
  not g15151 (n_7266, n8125);
  and g15152 (n8139, n_7266, n8138);
  not g15153 (n_7267, n8138);
  and g15154 (n8140, n8125, n_7267);
  not g15155 (n_7268, n8139);
  not g15156 (n_7269, n8140);
  and g15157 (n8141, n_7268, n_7269);
  not g15158 (n_7270, n8124);
  and g15159 (n8142, n_7270, n8141);
  not g15160 (n_7271, n8141);
  and g15161 (n8143, n8124, n_7271);
  not g15162 (n_7272, n8142);
  not g15163 (n_7273, n8143);
  and g15164 (n8144, n_7272, n_7273);
  not g15165 (n_7274, n8123);
  and g15166 (n8145, n_7274, n8144);
  not g15167 (n_7275, n8144);
  and g15168 (n8146, n8123, n_7275);
  not g15169 (n_7276, n8145);
  not g15170 (n_7277, n8146);
  and g15171 (n8147, n_7276, n_7277);
  not g15172 (n_7278, n8147);
  and g15173 (n8148, n8122, n_7278);
  not g15174 (n_7279, n8122);
  and g15175 (n8149, n_7279, n8147);
  not g15176 (n_7280, n8148);
  not g15177 (n_7281, n8149);
  and g15178 (n8150, n_7280, n_7281);
  and g15179 (n8151, n_7020, n_7024);
  and g15180 (n8152, n_7051, n_7056);
  and g15181 (n8153, n606, n5250);
  and g15182 (n8154, n602, n6252);
  and g15183 (n8155, \a[45] , \a[48] );
  and g15184 (n8156, n1605, n8155);
  not g15185 (n_7282, n8154);
  not g15186 (n_7283, n8156);
  and g15187 (n8157, n_7282, n_7283);
  not g15188 (n_7284, n8153);
  not g15189 (n_7285, n8157);
  and g15190 (n8158, n_7284, n_7285);
  not g15191 (n_7286, n8158);
  and g15192 (n8159, n_7284, n_7286);
  and g15193 (n8160, \a[12] , \a[47] );
  and g15194 (n8161, \a[14] , \a[45] );
  not g15195 (n_7287, n8160);
  not g15196 (n_7288, n8161);
  and g15197 (n8162, n_7287, n_7288);
  not g15198 (n_7289, n8162);
  and g15199 (n8163, n8159, n_7289);
  and g15200 (n8164, \a[48] , n_7286);
  and g15201 (n8165, \a[11] , n8164);
  not g15202 (n_7290, n8163);
  not g15203 (n_7291, n8165);
  and g15204 (n8166, n_7290, n_7291);
  and g15205 (n8167, \a[13] , \a[46] );
  and g15206 (n8168, \a[28] , \a[31] );
  not g15207 (n_7292, n2617);
  not g15208 (n_7293, n8168);
  and g15209 (n8169, n_7292, n_7293);
  and g15210 (n8170, n2617, n8168);
  not g15211 (n_7294, n8170);
  and g15212 (n8171, n8167, n_7294);
  not g15213 (n_7295, n8169);
  and g15214 (n8172, n_7295, n8171);
  not g15215 (n_7296, n8172);
  and g15216 (n8173, n8167, n_7296);
  and g15217 (n8174, n_7294, n_7296);
  and g15218 (n8175, n_7295, n8174);
  not g15219 (n_7297, n8173);
  not g15220 (n_7298, n8175);
  and g15221 (n8176, n_7297, n_7298);
  not g15222 (n_7299, n8166);
  not g15223 (n_7300, n8176);
  and g15224 (n8177, n_7299, n_7300);
  not g15225 (n_7301, n8177);
  and g15226 (n8178, n_7299, n_7301);
  and g15227 (n8179, n_7300, n_7301);
  not g15228 (n_7302, n8178);
  not g15229 (n_7303, n8179);
  and g15230 (n8180, n_7302, n_7303);
  and g15231 (n8181, \a[16] , \a[43] );
  and g15232 (n8182, \a[17] , \a[42] );
  not g15233 (n_7304, n8181);
  not g15234 (n_7305, n8182);
  and g15235 (n8183, n_7304, n_7305);
  and g15236 (n8184, n1048, n5018);
  not g15237 (n_7306, n8184);
  not g15240 (n_7307, n8183);
  not g15242 (n_7308, n8187);
  and g15243 (n8188, \a[51] , n_7308);
  and g15244 (n8189, \a[8] , n8188);
  and g15245 (n8190, n_7306, n_7308);
  and g15246 (n8191, n_7307, n8190);
  not g15247 (n_7309, n8189);
  not g15248 (n_7310, n8191);
  and g15249 (n8192, n_7309, n_7310);
  not g15250 (n_7311, n8180);
  not g15251 (n_7312, n8192);
  and g15252 (n8193, n_7311, n_7312);
  not g15253 (n_7313, n8193);
  and g15254 (n8194, n_7311, n_7313);
  and g15255 (n8195, n_7312, n_7313);
  not g15256 (n_7314, n8194);
  not g15257 (n_7315, n8195);
  and g15258 (n8196, n_7314, n_7315);
  and g15259 (n8197, \a[2] , \a[57] );
  and g15260 (n8198, \a[3] , \a[56] );
  not g15261 (n_7316, n8197);
  not g15262 (n_7317, n8198);
  and g15263 (n8199, n_7316, n_7317);
  and g15264 (n8200, \a[56] , \a[57] );
  and g15265 (n8201, n218, n8200);
  not g15266 (n_7318, n8199);
  not g15267 (n_7319, n8201);
  and g15268 (n8202, n_7318, n_7319);
  and g15269 (n8203, n7897, n8202);
  not g15270 (n_7320, n8203);
  and g15271 (n8204, n_7319, n_7320);
  and g15272 (n8205, n_7318, n8204);
  and g15273 (n8206, n7897, n_7320);
  not g15274 (n_7321, n8205);
  not g15275 (n_7322, n8206);
  and g15276 (n8207, n_7321, n_7322);
  not g15277 (n_7323, n8207);
  and g15278 (n8208, n8025, n_7323);
  not g15279 (n_7324, n8025);
  and g15280 (n8209, n_7324, n8207);
  not g15281 (n_7325, n8208);
  not g15282 (n_7326, n8209);
  and g15283 (n8210, n_7325, n_7326);
  and g15284 (n8211, n226, n7701);
  and g15285 (n8212, \a[19] , \a[55] );
  and g15286 (n8213, n4583, n8212);
  not g15287 (n_7327, n8211);
  not g15288 (n_7328, n8213);
  and g15289 (n8214, n_7327, n_7328);
  and g15290 (n8215, \a[5] , \a[54] );
  and g15291 (n8216, \a[19] , \a[40] );
  and g15292 (n8217, n8215, n8216);
  not g15293 (n_7329, n8214);
  not g15294 (n_7330, n8217);
  and g15295 (n8218, n_7329, n_7330);
  not g15296 (n_7331, n8218);
  and g15297 (n8219, \a[55] , n_7331);
  and g15298 (n8220, \a[4] , n8219);
  and g15299 (n8221, n_7330, n_7331);
  not g15300 (n_7332, n8215);
  not g15301 (n_7333, n8216);
  and g15302 (n8222, n_7332, n_7333);
  not g15303 (n_7334, n8222);
  and g15304 (n8223, n8221, n_7334);
  not g15305 (n_7335, n8220);
  not g15306 (n_7336, n8223);
  and g15307 (n8224, n_7335, n_7336);
  not g15308 (n_7337, n8210);
  not g15309 (n_7338, n8224);
  and g15310 (n8225, n_7337, n_7338);
  and g15311 (n8226, n8210, n8224);
  not g15312 (n_7339, n8225);
  not g15313 (n_7340, n8226);
  and g15314 (n8227, n_7339, n_7340);
  not g15315 (n_7341, n8227);
  and g15316 (n8228, n8196, n_7341);
  not g15317 (n_7342, n8196);
  and g15318 (n8229, n_7342, n8227);
  not g15319 (n_7343, n8228);
  not g15320 (n_7344, n8229);
  and g15321 (n8230, n_7343, n_7344);
  not g15322 (n_7345, n8152);
  and g15323 (n8231, n_7345, n8230);
  not g15324 (n_7346, n8230);
  and g15325 (n8232, n8152, n_7346);
  not g15326 (n_7347, n8231);
  not g15327 (n_7348, n8232);
  and g15328 (n8233, n_7347, n_7348);
  not g15329 (n_7349, n8233);
  and g15330 (n8234, n8151, n_7349);
  not g15331 (n_7350, n8151);
  and g15332 (n8235, n_7350, n8233);
  not g15333 (n_7351, n8234);
  not g15334 (n_7352, n8235);
  and g15335 (n8236, n_7351, n_7352);
  and g15336 (n8237, \a[18] , \a[52] );
  and g15337 (n8238, n5411, n8237);
  and g15338 (n8239, \a[41] , \a[53] );
  and g15339 (n8240, n1478, n8239);
  and g15340 (n8241, n335, n7433);
  not g15341 (n_7353, n8240);
  not g15342 (n_7354, n8241);
  and g15343 (n8242, n_7353, n_7354);
  not g15344 (n_7355, n8238);
  not g15345 (n_7356, n8242);
  and g15346 (n8243, n_7355, n_7356);
  not g15347 (n_7357, n8243);
  and g15348 (n8244, n_7355, n_7357);
  and g15349 (n8245, \a[7] , \a[52] );
  and g15350 (n8246, \a[18] , \a[41] );
  not g15351 (n_7358, n8245);
  not g15352 (n_7359, n8246);
  and g15353 (n8247, n_7358, n_7359);
  not g15354 (n_7360, n8247);
  and g15355 (n8248, n8244, n_7360);
  and g15356 (n8249, \a[53] , n_7357);
  and g15357 (n8250, \a[6] , n8249);
  not g15358 (n_7361, n8248);
  not g15359 (n_7362, n8250);
  and g15360 (n8251, n_7361, n_7362);
  and g15361 (n8252, \a[44] , \a[49] );
  and g15362 (n8253, n685, n8252);
  and g15363 (n8254, \a[44] , \a[50] );
  and g15364 (n8255, n1517, n8254);
  and g15365 (n8256, n484, n6325);
  not g15366 (n_7363, n8255);
  not g15367 (n_7364, n8256);
  and g15368 (n8257, n_7363, n_7364);
  not g15369 (n_7365, n8253);
  not g15370 (n_7366, n8257);
  and g15371 (n8258, n_7365, n_7366);
  not g15372 (n_7367, n8258);
  and g15373 (n8259, \a[50] , n_7367);
  and g15374 (n8260, \a[9] , n8259);
  and g15375 (n8261, \a[10] , \a[49] );
  not g15376 (n_7368, n5298);
  not g15377 (n_7369, n8261);
  and g15378 (n8262, n_7368, n_7369);
  and g15379 (n8263, n_7365, n_7367);
  not g15380 (n_7370, n8262);
  and g15381 (n8264, n_7370, n8263);
  not g15382 (n_7371, n8260);
  not g15383 (n_7372, n8264);
  and g15384 (n8265, n_7371, n_7372);
  not g15385 (n_7373, n8251);
  not g15386 (n_7374, n8265);
  and g15387 (n8266, n_7373, n_7374);
  not g15388 (n_7375, n8266);
  and g15389 (n8267, n_7373, n_7375);
  and g15390 (n8268, n_7374, n_7375);
  not g15391 (n_7376, n8267);
  not g15392 (n_7377, n8268);
  and g15393 (n8269, n_7376, n_7377);
  and g15394 (n8270, n_7045, n_7048);
  and g15395 (n8271, n8269, n8270);
  not g15396 (n_7378, n8269);
  not g15397 (n_7379, n8270);
  and g15398 (n8272, n_7378, n_7379);
  not g15399 (n_7380, n8271);
  not g15400 (n_7381, n8272);
  and g15401 (n8273, n_7380, n_7381);
  and g15402 (n8274, n_7013, n_7017);
  not g15403 (n_7382, n8273);
  and g15404 (n8275, n_7382, n8274);
  not g15405 (n_7383, n8274);
  and g15406 (n8276, n8273, n_7383);
  not g15407 (n_7384, n8275);
  not g15408 (n_7385, n8276);
  and g15409 (n8277, n_7384, n_7385);
  and g15410 (n8278, n1574, n4565);
  and g15411 (n8279, n1693, n5430);
  and g15412 (n8280, n1494, n5083);
  not g15413 (n_7386, n8279);
  not g15414 (n_7387, n8280);
  and g15415 (n8281, n_7386, n_7387);
  not g15416 (n_7388, n8278);
  not g15417 (n_7389, n8281);
  and g15418 (n8282, n_7388, n_7389);
  not g15419 (n_7390, n8282);
  and g15420 (n8283, n_7388, n_7390);
  and g15421 (n8284, \a[21] , \a[38] );
  and g15422 (n8285, \a[22] , \a[37] );
  not g15423 (n_7391, n8284);
  not g15424 (n_7392, n8285);
  and g15425 (n8286, n_7391, n_7392);
  not g15426 (n_7393, n8286);
  and g15427 (n8287, n8283, n_7393);
  and g15428 (n8288, \a[39] , n_7390);
  and g15429 (n8289, \a[20] , n8288);
  not g15430 (n_7394, n8287);
  not g15431 (n_7395, n8289);
  and g15432 (n8290, n_7394, n_7395);
  and g15433 (n8291, n1904, n3319);
  and g15434 (n8292, n1547, n4595);
  and g15435 (n8293, n1666, n3828);
  not g15436 (n_7396, n8292);
  not g15437 (n_7397, n8293);
  and g15438 (n8294, n_7396, n_7397);
  not g15439 (n_7398, n8291);
  not g15440 (n_7399, n8294);
  and g15441 (n8295, n_7398, n_7399);
  not g15442 (n_7400, n8295);
  and g15443 (n8296, \a[36] , n_7400);
  and g15444 (n8297, \a[23] , n8296);
  and g15445 (n8298, \a[24] , \a[35] );
  and g15446 (n8299, \a[25] , \a[34] );
  not g15447 (n_7401, n8298);
  not g15448 (n_7402, n8299);
  and g15449 (n8300, n_7401, n_7402);
  and g15450 (n8301, n_7398, n_7400);
  not g15451 (n_7403, n8300);
  and g15452 (n8302, n_7403, n8301);
  not g15453 (n_7404, n8297);
  not g15454 (n_7405, n8302);
  and g15455 (n8303, n_7404, n_7405);
  not g15456 (n_7406, n8290);
  not g15457 (n_7407, n8303);
  and g15458 (n8304, n_7406, n_7407);
  not g15459 (n_7408, n8304);
  and g15460 (n8305, n_7406, n_7408);
  and g15461 (n8306, n_7407, n_7408);
  not g15462 (n_7409, n8305);
  not g15463 (n_7410, n8306);
  and g15464 (n8307, n_7409, n_7410);
  and g15465 (n8308, \a[32] , \a[59] );
  and g15466 (n8309, n1812, n8308);
  and g15467 (n8310, n2227, n3143);
  and g15468 (n8311, \a[26] , \a[59] );
  and g15469 (n8312, n2605, n8311);
  not g15470 (n_7412, n8310);
  not g15471 (n_7413, n8312);
  and g15472 (n8313, n_7412, n_7413);
  not g15473 (n_7414, n8309);
  not g15474 (n_7415, n8313);
  and g15475 (n8314, n_7414, n_7415);
  not g15476 (n_7416, n8314);
  and g15477 (n8315, \a[33] , n_7416);
  and g15478 (n8316, \a[26] , n8315);
  and g15479 (n8317, n_7414, n_7416);
  and g15480 (n8318, \a[0] , \a[59] );
  and g15481 (n8319, \a[27] , \a[32] );
  not g15482 (n_7417, n8318);
  not g15483 (n_7418, n8319);
  and g15484 (n8320, n_7417, n_7418);
  not g15485 (n_7419, n8320);
  and g15486 (n8321, n8317, n_7419);
  not g15487 (n_7420, n8316);
  not g15488 (n_7421, n8321);
  and g15489 (n8322, n_7420, n_7421);
  not g15490 (n_7422, n8307);
  not g15491 (n_7423, n8322);
  and g15492 (n8323, n_7422, n_7423);
  not g15493 (n_7424, n8323);
  and g15494 (n8324, n_7422, n_7424);
  and g15495 (n8325, n_7423, n_7424);
  not g15496 (n_7425, n8324);
  not g15497 (n_7426, n8325);
  and g15498 (n8326, n_7425, n_7426);
  not g15499 (n_7427, n8326);
  and g15500 (n8327, n8277, n_7427);
  not g15501 (n_7428, n8277);
  and g15502 (n8328, n_7428, n8326);
  not g15503 (n_7429, n8328);
  and g15504 (n8329, n8236, n_7429);
  not g15505 (n_7430, n8327);
  and g15506 (n8330, n_7430, n8329);
  not g15507 (n_7431, n8330);
  and g15508 (n8331, n8236, n_7431);
  and g15509 (n8332, n_7429, n_7431);
  and g15510 (n8333, n_7430, n8332);
  not g15511 (n_7432, n8331);
  not g15512 (n_7433, n8333);
  and g15513 (n8334, n_7432, n_7433);
  and g15514 (n8335, n_7029, n_7033);
  and g15515 (n8336, n_7211, n_7223);
  and g15516 (n8337, n_7151, n_7166);
  and g15517 (n8338, n8336, n8337);
  not g15518 (n_7434, n8336);
  not g15519 (n_7435, n8337);
  and g15520 (n8339, n_7434, n_7435);
  not g15521 (n_7436, n8338);
  not g15522 (n_7437, n8339);
  and g15523 (n8340, n_7436, n_7437);
  and g15524 (n8341, n_7114, n_7129);
  not g15525 (n_7438, n8340);
  and g15526 (n8342, n_7438, n8341);
  not g15527 (n_7439, n8341);
  and g15528 (n8343, n8340, n_7439);
  not g15529 (n_7440, n8342);
  not g15530 (n_7441, n8343);
  and g15531 (n8344, n_7440, n_7441);
  and g15532 (n8345, n_7169, n_7170);
  not g15533 (n_7442, n8345);
  and g15534 (n8346, n_7176, n_7442);
  and g15535 (n8347, n7950, n8090);
  not g15536 (n_7443, n7950);
  not g15537 (n_7444, n8090);
  and g15538 (n8348, n_7443, n_7444);
  not g15539 (n_7445, n8347);
  not g15540 (n_7446, n8348);
  and g15541 (n8349, n_7445, n_7446);
  not g15542 (n_7447, n8349);
  and g15543 (n8350, n7983, n_7447);
  not g15544 (n_7448, n7983);
  and g15545 (n8351, n_7448, n8349);
  not g15546 (n_7449, n8350);
  not g15547 (n_7450, n8351);
  and g15548 (n8352, n_7449, n_7450);
  and g15549 (n8353, n7965, n8009);
  not g15550 (n_7451, n7965);
  not g15551 (n_7452, n8009);
  and g15552 (n8354, n_7451, n_7452);
  not g15553 (n_7453, n8353);
  not g15554 (n_7454, n8354);
  and g15555 (n8355, n_7453, n_7454);
  not g15556 (n_7455, n8355);
  and g15557 (n8356, n7997, n_7455);
  not g15558 (n_7456, n7997);
  and g15559 (n8357, n_7456, n8355);
  not g15560 (n_7457, n8356);
  not g15561 (n_7458, n8357);
  and g15562 (n8358, n_7457, n_7458);
  and g15563 (n8359, \a[58] , n2402);
  and g15564 (n8360, \a[1] , \a[58] );
  not g15565 (n_7459, \a[30] );
  not g15566 (n_7460, n8360);
  and g15567 (n8361, n_7459, n_7460);
  not g15568 (n_7461, n8359);
  not g15569 (n_7462, n8361);
  and g15570 (n8362, n_7461, n_7462);
  not g15571 (n_7463, n8362);
  and g15572 (n8363, n8072, n_7463);
  not g15573 (n_7464, n8072);
  and g15574 (n8364, n_7464, n8362);
  not g15575 (n_7465, n8363);
  not g15576 (n_7466, n8364);
  and g15577 (n8365, n_7465, n_7466);
  not g15578 (n_7467, n8059);
  and g15579 (n8366, n_7467, n8365);
  not g15580 (n_7468, n8365);
  and g15581 (n8367, n8059, n_7468);
  not g15582 (n_7469, n8366);
  not g15583 (n_7470, n8367);
  and g15584 (n8368, n_7469, n_7470);
  and g15585 (n8369, n8358, n8368);
  not g15586 (n_7471, n8369);
  and g15587 (n8370, n8358, n_7471);
  and g15588 (n8371, n8368, n_7471);
  not g15589 (n_7472, n8370);
  not g15590 (n_7473, n8371);
  and g15591 (n8372, n_7472, n_7473);
  not g15592 (n_7474, n8372);
  and g15593 (n8373, n8352, n_7474);
  not g15594 (n_7475, n8352);
  and g15595 (n8374, n_7475, n_7473);
  and g15596 (n8375, n_7472, n8374);
  not g15597 (n_7476, n8373);
  not g15598 (n_7477, n8375);
  and g15599 (n8376, n_7476, n_7477);
  not g15600 (n_7478, n8346);
  and g15601 (n8377, n_7478, n8376);
  not g15602 (n_7479, n8377);
  and g15603 (n8378, n_7478, n_7479);
  and g15604 (n8379, n8376, n_7479);
  not g15605 (n_7480, n8378);
  not g15606 (n_7481, n8379);
  and g15607 (n8380, n_7480, n_7481);
  not g15608 (n_7482, n8380);
  and g15609 (n8381, n8344, n_7482);
  not g15610 (n_7483, n8344);
  and g15611 (n8382, n_7483, n_7481);
  and g15612 (n8383, n_7480, n8382);
  not g15613 (n_7484, n8381);
  not g15614 (n_7485, n8383);
  and g15615 (n8384, n_7484, n_7485);
  not g15616 (n_7486, n8335);
  and g15617 (n8385, n_7486, n8384);
  not g15618 (n_7487, n8384);
  and g15619 (n8386, n8335, n_7487);
  not g15620 (n_7488, n8385);
  not g15621 (n_7489, n8386);
  and g15622 (n8387, n_7488, n_7489);
  not g15623 (n_7490, n8334);
  and g15624 (n8388, n_7490, n8387);
  not g15625 (n_7491, n8387);
  and g15626 (n8389, n8334, n_7491);
  not g15627 (n_7492, n8388);
  not g15628 (n_7493, n8389);
  and g15629 (n8390, n_7492, n_7493);
  and g15630 (n8391, n8150, n8390);
  not g15631 (n_7494, n8150);
  not g15632 (n_7495, n8390);
  and g15633 (n8392, n_7494, n_7495);
  not g15634 (n_7496, n8391);
  not g15635 (n_7497, n8392);
  and g15636 (n8393, n_7496, n_7497);
  and g15637 (n8394, n_7038, n_7245);
  not g15638 (n_7498, n8393);
  and g15639 (n8395, n_7498, n8394);
  not g15640 (n_7499, n8394);
  and g15641 (n8396, n8393, n_7499);
  not g15642 (n_7500, n8395);
  not g15643 (n_7501, n8396);
  and g15644 (n8397, n_7500, n_7501);
  not g15645 (n_7502, n8119);
  and g15646 (n8398, n_7248, n_7502);
  not g15647 (n_7503, n8397);
  and g15648 (n8399, n_7503, n8398);
  not g15649 (n_7504, n8398);
  and g15650 (n8400, n8397, n_7504);
  not g15651 (n_7505, n8399);
  not g15652 (n_7506, n8400);
  and g15653 (\asquared[60] , n_7505, n_7506);
  and g15654 (n8402, n_7281, n_7496);
  and g15655 (n8403, n_7488, n_7492);
  and g15656 (n8404, n_7352, n_7431);
  and g15657 (n8405, n_7479, n_7484);
  and g15658 (n8406, n_7454, n_7458);
  and g15659 (n8407, n_7446, n_7450);
  and g15660 (n8408, n8406, n8407);
  not g15661 (n_7507, n8406);
  not g15662 (n_7508, n8407);
  and g15663 (n8409, n_7507, n_7508);
  not g15664 (n_7509, n8408);
  not g15665 (n_7510, n8409);
  and g15666 (n8410, n_7509, n_7510);
  and g15667 (n8411, n_7324, n_7323);
  not g15668 (n_7511, n8411);
  and g15669 (n8412, n_7339, n_7511);
  not g15670 (n_7512, n8410);
  and g15671 (n8413, n_7512, n8412);
  not g15672 (n_7513, n8412);
  and g15673 (n8414, n8410, n_7513);
  not g15674 (n_7514, n8413);
  not g15675 (n_7515, n8414);
  and g15676 (n8415, n_7514, n_7515);
  and g15677 (n8416, n_7437, n_7441);
  not g15678 (n_7516, n8415);
  and g15679 (n8417, n_7516, n8416);
  not g15680 (n_7517, n8416);
  and g15681 (n8418, n8415, n_7517);
  not g15682 (n_7518, n8417);
  not g15683 (n_7519, n8418);
  and g15684 (n8419, n_7518, n_7519);
  and g15685 (n8420, n_7385, n_7430);
  not g15686 (n_7520, n8420);
  and g15687 (n8421, n8419, n_7520);
  not g15688 (n_7521, n8419);
  and g15689 (n8422, n_7521, n8420);
  not g15690 (n_7522, n8421);
  not g15691 (n_7523, n8422);
  and g15692 (n8423, n_7522, n_7523);
  not g15693 (n_7524, n8405);
  and g15694 (n8424, n_7524, n8423);
  not g15695 (n_7525, n8423);
  and g15696 (n8425, n8405, n_7525);
  not g15697 (n_7526, n8424);
  not g15698 (n_7527, n8425);
  and g15699 (n8426, n_7526, n_7527);
  not g15700 (n_7528, n8404);
  and g15701 (n8427, n_7528, n8426);
  not g15702 (n_7529, n8426);
  and g15703 (n8428, n8404, n_7529);
  not g15704 (n_7530, n8427);
  not g15705 (n_7531, n8428);
  and g15706 (n8429, n_7530, n_7531);
  not g15707 (n_7532, n8429);
  and g15708 (n8430, n8403, n_7532);
  not g15709 (n_7533, n8403);
  and g15710 (n8431, n_7533, n8429);
  not g15711 (n_7534, n8430);
  not g15712 (n_7535, n8431);
  and g15713 (n8432, n_7534, n_7535);
  and g15714 (n8433, n_7264, n_7268);
  and g15715 (n8434, n209, n8200);
  and g15716 (n8435, n252, n7942);
  and g15717 (n8436, \a[57] , \a[58] );
  and g15718 (n8437, n218, n8436);
  not g15719 (n_7536, n8435);
  not g15720 (n_7537, n8437);
  and g15721 (n8438, n_7536, n_7537);
  not g15722 (n_7538, n8434);
  not g15723 (n_7539, n8438);
  and g15724 (n8439, n_7538, n_7539);
  not g15725 (n_7540, n8439);
  and g15726 (n8440, n_7538, n_7540);
  and g15727 (n8441, \a[3] , \a[57] );
  and g15728 (n8442, \a[4] , \a[56] );
  not g15729 (n_7541, n8441);
  not g15730 (n_7542, n8442);
  and g15731 (n8443, n_7541, n_7542);
  not g15732 (n_7543, n8443);
  and g15733 (n8444, n8440, n_7543);
  and g15734 (n8445, \a[58] , n_7540);
  and g15735 (n8446, \a[2] , n8445);
  not g15736 (n_7544, n8444);
  not g15737 (n_7545, n8446);
  and g15738 (n8447, n_7544, n_7545);
  and g15739 (n8448, n1574, n5083);
  and g15740 (n8449, n1693, n3803);
  and g15741 (n8450, n1494, n4171);
  not g15742 (n_7546, n8449);
  not g15743 (n_7547, n8450);
  and g15744 (n8451, n_7546, n_7547);
  not g15745 (n_7548, n8448);
  not g15746 (n_7549, n8451);
  and g15747 (n8452, n_7548, n_7549);
  not g15748 (n_7550, n8452);
  and g15749 (n8453, \a[40] , n_7550);
  and g15750 (n8454, \a[20] , n8453);
  and g15751 (n8455, \a[21] , \a[39] );
  and g15752 (n8456, \a[22] , \a[38] );
  not g15753 (n_7551, n8455);
  not g15754 (n_7552, n8456);
  and g15755 (n8457, n_7551, n_7552);
  and g15756 (n8458, n_7548, n_7550);
  not g15757 (n_7553, n8457);
  and g15758 (n8459, n_7553, n8458);
  not g15759 (n_7554, n8454);
  not g15760 (n_7555, n8459);
  and g15761 (n8460, n_7554, n_7555);
  not g15762 (n_7556, n8447);
  not g15763 (n_7557, n8460);
  and g15764 (n8461, n_7556, n_7557);
  not g15765 (n_7558, n8461);
  and g15766 (n8462, n_7556, n_7558);
  and g15767 (n8463, n_7557, n_7558);
  not g15768 (n_7559, n8462);
  not g15769 (n_7560, n8463);
  and g15770 (n8464, n_7559, n_7560);
  and g15771 (n8465, n2463, n3319);
  and g15772 (n8466, n2301, n4595);
  and g15773 (n8467, n1904, n3828);
  not g15774 (n_7561, n8466);
  not g15775 (n_7562, n8467);
  and g15776 (n8468, n_7561, n_7562);
  not g15777 (n_7563, n8465);
  not g15778 (n_7564, n8468);
  and g15779 (n8469, n_7563, n_7564);
  not g15780 (n_7565, n8469);
  and g15781 (n8470, \a[36] , n_7565);
  and g15782 (n8471, \a[24] , n8470);
  and g15783 (n8472, n_7563, n_7565);
  and g15784 (n8473, \a[25] , \a[35] );
  and g15785 (n8474, \a[26] , \a[34] );
  not g15786 (n_7566, n8473);
  not g15787 (n_7567, n8474);
  and g15788 (n8475, n_7566, n_7567);
  not g15789 (n_7568, n8475);
  and g15790 (n8476, n8472, n_7568);
  not g15791 (n_7569, n8471);
  not g15792 (n_7570, n8476);
  and g15793 (n8477, n_7569, n_7570);
  not g15794 (n_7571, n8464);
  not g15795 (n_7572, n8477);
  and g15796 (n8478, n_7571, n_7572);
  not g15797 (n_7573, n8478);
  and g15798 (n8479, n_7571, n_7573);
  and g15799 (n8480, n_7572, n_7573);
  not g15800 (n_7574, n8479);
  not g15801 (n_7575, n8480);
  and g15802 (n8481, n_7574, n_7575);
  and g15803 (n8482, n_7257, n_7261);
  and g15804 (n8483, n8481, n8482);
  not g15805 (n_7576, n8481);
  not g15806 (n_7577, n8482);
  and g15807 (n8484, n_7576, n_7577);
  not g15808 (n_7578, n8483);
  not g15809 (n_7579, n8484);
  and g15810 (n8485, n_7578, n_7579);
  and g15811 (n8486, \a[44] , \a[51] );
  and g15812 (n8487, n847, n8486);
  and g15813 (n8488, n1048, n5296);
  and g15814 (n8489, n6516, n7772);
  not g15815 (n_7580, n8488);
  not g15816 (n_7581, n8489);
  and g15817 (n8490, n_7580, n_7581);
  not g15818 (n_7582, n8487);
  not g15819 (n_7583, n8490);
  and g15820 (n8491, n_7582, n_7583);
  not g15821 (n_7584, n8491);
  and g15822 (n8492, \a[43] , n_7584);
  and g15823 (n8493, \a[17] , n8492);
  and g15824 (n8494, n_7582, n_7584);
  and g15825 (n8495, \a[9] , \a[51] );
  and g15826 (n8496, \a[16] , \a[44] );
  not g15827 (n_7585, n8495);
  not g15828 (n_7586, n8496);
  and g15829 (n8497, n_7585, n_7586);
  not g15830 (n_7587, n8497);
  and g15831 (n8498, n8494, n_7587);
  not g15832 (n_7588, n8493);
  not g15833 (n_7589, n8498);
  and g15834 (n8499, n_7588, n_7589);
  not g15835 (n_7590, n8499);
  and g15836 (n8500, n8159, n_7590);
  not g15837 (n_7591, n8159);
  and g15838 (n8501, n_7591, n8499);
  not g15839 (n_7592, n8500);
  not g15840 (n_7593, n8501);
  and g15841 (n8502, n_7592, n_7593);
  and g15842 (n8503, \a[45] , \a[49] );
  and g15843 (n8504, n816, n8503);
  and g15844 (n8505, n723, n6325);
  and g15845 (n8506, \a[45] , \a[50] );
  and g15846 (n8507, n685, n8506);
  not g15847 (n_7594, n8505);
  not g15848 (n_7595, n8507);
  and g15849 (n8508, n_7594, n_7595);
  not g15850 (n_7596, n8504);
  not g15851 (n_7597, n8508);
  and g15852 (n8509, n_7596, n_7597);
  not g15853 (n_7598, n8509);
  and g15854 (n8510, \a[50] , n_7598);
  and g15855 (n8511, \a[10] , n8510);
  and g15856 (n8512, \a[11] , \a[49] );
  and g15857 (n8513, \a[15] , \a[45] );
  not g15858 (n_7599, n8512);
  not g15859 (n_7600, n8513);
  and g15860 (n8514, n_7599, n_7600);
  and g15861 (n8515, n_7596, n_7598);
  not g15862 (n_7601, n8514);
  and g15863 (n8516, n_7601, n8515);
  not g15864 (n_7602, n8511);
  not g15865 (n_7603, n8516);
  and g15866 (n8517, n_7602, n_7603);
  not g15867 (n_7604, n8502);
  not g15868 (n_7605, n8517);
  and g15869 (n8518, n_7604, n_7605);
  and g15870 (n8519, n8502, n8517);
  not g15871 (n_7606, n8518);
  not g15872 (n_7607, n8519);
  and g15873 (n8520, n_7606, n_7607);
  not g15874 (n_7608, n8485);
  not g15875 (n_7609, n8520);
  and g15876 (n8521, n_7608, n_7609);
  and g15877 (n8522, n8485, n8520);
  not g15878 (n_7610, n8521);
  not g15879 (n_7611, n8522);
  and g15880 (n8523, n_7610, n_7611);
  not g15881 (n_7612, n8433);
  and g15882 (n8524, n_7612, n8523);
  not g15883 (n_7613, n8524);
  and g15884 (n8525, n_7612, n_7613);
  and g15885 (n8526, n8523, n_7613);
  not g15886 (n_7614, n8525);
  not g15887 (n_7615, n8526);
  and g15888 (n8527, n_7614, n_7615);
  and g15889 (n8528, n_7471, n_7476);
  and g15890 (n8529, \a[0] , \a[60] );
  and g15891 (n8530, n8359, n8529);
  not g15892 (n_7617, n8530);
  and g15893 (n8531, n8359, n_7617);
  and g15894 (n8532, n_7461, n8529);
  not g15895 (n_7618, n8531);
  not g15896 (n_7619, n8532);
  and g15897 (n8533, n_7618, n_7619);
  and g15898 (n8534, \a[1] , \a[59] );
  and g15899 (n8535, n3452, n8534);
  not g15900 (n_7620, n8535);
  and g15901 (n8536, n8534, n_7620);
  and g15902 (n8537, n3452, n_7620);
  not g15903 (n_7621, n8536);
  not g15904 (n_7622, n8537);
  and g15905 (n8538, n_7621, n_7622);
  not g15906 (n_7623, n8533);
  not g15907 (n_7624, n8538);
  and g15908 (n8539, n_7623, n_7624);
  not g15909 (n_7625, n8539);
  and g15910 (n8540, n_7623, n_7625);
  and g15911 (n8541, n_7624, n_7625);
  not g15912 (n_7626, n8540);
  not g15913 (n_7627, n8541);
  and g15914 (n8542, n_7626, n_7627);
  and g15915 (n8543, n2331, n3143);
  and g15916 (n8544, n4059, n7377);
  not g15917 (n_7628, n8543);
  not g15918 (n_7629, n8544);
  and g15919 (n8545, n_7628, n_7629);
  and g15920 (n8546, \a[23] , \a[37] );
  and g15921 (n8547, n5863, n8546);
  not g15922 (n_7630, n8545);
  not g15923 (n_7631, n8547);
  and g15924 (n8548, n_7630, n_7631);
  not g15925 (n_7632, n8548);
  and g15926 (n8549, \a[33] , n_7632);
  and g15927 (n8550, \a[27] , n8549);
  and g15928 (n8551, n_7631, n_7632);
  not g15929 (n_7633, n5863);
  not g15930 (n_7634, n8546);
  and g15931 (n8552, n_7633, n_7634);
  not g15932 (n_7635, n8552);
  and g15933 (n8553, n8551, n_7635);
  not g15934 (n_7636, n8550);
  not g15935 (n_7637, n8553);
  and g15936 (n8554, n_7636, n_7637);
  not g15937 (n_7638, n8542);
  not g15938 (n_7639, n8554);
  and g15939 (n8555, n_7638, n_7639);
  not g15940 (n_7640, n8555);
  and g15941 (n8556, n_7638, n_7640);
  and g15942 (n8557, n_7639, n_7640);
  not g15943 (n_7641, n8556);
  not g15944 (n_7642, n8557);
  and g15945 (n8558, n_7641, n_7642);
  and g15946 (n8559, n_7466, n_7469);
  and g15947 (n8560, n8558, n8559);
  not g15948 (n_7643, n8558);
  not g15949 (n_7644, n8559);
  and g15950 (n8561, n_7643, n_7644);
  not g15951 (n_7645, n8560);
  not g15952 (n_7646, n8561);
  and g15953 (n8562, n_7645, n_7646);
  and g15954 (n8563, n380, n7433);
  and g15955 (n8564, \a[18] , \a[53] );
  and g15956 (n8565, n5619, n8564);
  not g15957 (n_7647, n8563);
  not g15958 (n_7648, n8565);
  and g15959 (n8566, n_7647, n_7648);
  and g15960 (n8567, \a[8] , \a[52] );
  and g15961 (n8568, \a[18] , \a[42] );
  and g15962 (n8569, n8567, n8568);
  not g15963 (n_7649, n8566);
  not g15964 (n_7650, n8569);
  and g15965 (n8570, n_7649, n_7650);
  not g15966 (n_7651, n8570);
  and g15967 (n8571, n_7650, n_7651);
  not g15968 (n_7652, n8567);
  not g15969 (n_7653, n8568);
  and g15970 (n8572, n_7652, n_7653);
  not g15971 (n_7654, n8572);
  and g15972 (n8573, n8571, n_7654);
  and g15973 (n8574, \a[53] , n_7651);
  and g15974 (n8575, \a[7] , n8574);
  not g15975 (n_7655, n8573);
  not g15976 (n_7656, n8575);
  and g15977 (n8576, n_7655, n_7656);
  and g15978 (n8577, n748, n6252);
  and g15979 (n8578, \a[46] , \a[48] );
  and g15980 (n8579, n606, n8578);
  and g15981 (n8580, n745, n5666);
  not g15982 (n_7657, n8579);
  not g15983 (n_7658, n8580);
  and g15984 (n8581, n_7657, n_7658);
  not g15985 (n_7659, n8577);
  not g15986 (n_7660, n8581);
  and g15987 (n8582, n_7659, n_7660);
  not g15988 (n_7661, n8582);
  and g15989 (n8583, n7400, n_7661);
  and g15990 (n8584, n_7659, n_7661);
  and g15991 (n8585, \a[12] , \a[48] );
  and g15992 (n8586, \a[13] , \a[47] );
  not g15993 (n_7662, n8585);
  not g15994 (n_7663, n8586);
  and g15995 (n8587, n_7662, n_7663);
  not g15996 (n_7664, n8587);
  and g15997 (n8588, n8584, n_7664);
  not g15998 (n_7665, n8583);
  not g15999 (n_7666, n8588);
  and g16000 (n8589, n_7665, n_7666);
  not g16001 (n_7667, n8576);
  not g16002 (n_7668, n8589);
  and g16003 (n8590, n_7667, n_7668);
  not g16004 (n_7669, n8590);
  and g16005 (n8591, n_7667, n_7669);
  and g16006 (n8592, n_7668, n_7669);
  not g16007 (n_7670, n8591);
  not g16008 (n_7671, n8592);
  and g16009 (n8593, n_7670, n_7671);
  and g16010 (n8594, \a[41] , \a[55] );
  and g16011 (n8595, n1502, n8594);
  and g16012 (n8596, n332, n7701);
  not g16013 (n_7672, n8595);
  not g16014 (n_7673, n8596);
  and g16015 (n8597, n_7672, n_7673);
  and g16016 (n8598, \a[6] , \a[54] );
  and g16017 (n8599, \a[19] , \a[41] );
  and g16018 (n8600, n8598, n8599);
  not g16019 (n_7674, n8597);
  not g16020 (n_7675, n8600);
  and g16021 (n8601, n_7674, n_7675);
  not g16022 (n_7676, n8601);
  and g16023 (n8602, \a[55] , n_7676);
  and g16024 (n8603, \a[5] , n8602);
  and g16025 (n8604, n_7675, n_7676);
  not g16026 (n_7677, n8598);
  not g16027 (n_7678, n8599);
  and g16028 (n8605, n_7677, n_7678);
  not g16029 (n_7679, n8605);
  and g16030 (n8606, n8604, n_7679);
  not g16031 (n_7680, n8603);
  not g16032 (n_7681, n8606);
  and g16033 (n8607, n_7680, n_7681);
  not g16034 (n_7682, n8593);
  not g16035 (n_7683, n8607);
  and g16036 (n8608, n_7682, n_7683);
  not g16037 (n_7684, n8608);
  and g16038 (n8609, n_7682, n_7684);
  and g16039 (n8610, n_7683, n_7684);
  not g16040 (n_7685, n8609);
  not g16041 (n_7686, n8610);
  and g16042 (n8611, n_7685, n_7686);
  not g16043 (n_7687, n8562);
  and g16044 (n8612, n_7687, n8611);
  not g16045 (n_7688, n8611);
  and g16046 (n8613, n8562, n_7688);
  not g16047 (n_7689, n8612);
  not g16048 (n_7690, n8613);
  and g16049 (n8614, n_7689, n_7690);
  not g16050 (n_7691, n8528);
  and g16051 (n8615, n_7691, n8614);
  not g16052 (n_7692, n8614);
  and g16053 (n8616, n8528, n_7692);
  not g16054 (n_7693, n8615);
  not g16055 (n_7694, n8616);
  and g16056 (n8617, n_7693, n_7694);
  not g16057 (n_7695, n8527);
  and g16058 (n8618, n_7695, n8617);
  not g16059 (n_7696, n8618);
  and g16060 (n8619, n8617, n_7696);
  and g16061 (n8620, n_7695, n_7696);
  not g16062 (n_7697, n8619);
  not g16063 (n_7698, n8620);
  and g16064 (n8621, n_7697, n_7698);
  and g16065 (n8622, n_7272, n_7276);
  and g16066 (n8623, n8190, n8244);
  not g16067 (n_7699, n8190);
  not g16068 (n_7700, n8244);
  and g16069 (n8624, n_7699, n_7700);
  not g16070 (n_7701, n8623);
  not g16071 (n_7702, n8624);
  and g16072 (n8625, n_7701, n_7702);
  not g16073 (n_7703, n8625);
  and g16074 (n8626, n8174, n_7703);
  not g16075 (n_7704, n8174);
  and g16076 (n8627, n_7704, n8625);
  not g16077 (n_7705, n8626);
  not g16078 (n_7706, n8627);
  and g16079 (n8628, n_7705, n_7706);
  and g16080 (n8629, n_7408, n_7424);
  not g16081 (n_7707, n8628);
  and g16082 (n8630, n_7707, n8629);
  not g16083 (n_7708, n8629);
  and g16084 (n8631, n8628, n_7708);
  not g16085 (n_7709, n8630);
  not g16086 (n_7710, n8631);
  and g16087 (n8632, n_7709, n_7710);
  and g16088 (n8633, n_7301, n_7313);
  not g16089 (n_7711, n8632);
  and g16090 (n8634, n_7711, n8633);
  not g16091 (n_7712, n8633);
  and g16092 (n8635, n8632, n_7712);
  not g16093 (n_7713, n8634);
  not g16094 (n_7714, n8635);
  and g16095 (n8636, n_7713, n_7714);
  and g16096 (n8637, n_7344, n_7347);
  and g16097 (n8638, n_7375, n_7381);
  and g16098 (n8639, n8221, n8283);
  not g16099 (n_7715, n8221);
  not g16100 (n_7716, n8283);
  and g16101 (n8640, n_7715, n_7716);
  not g16102 (n_7717, n8639);
  not g16103 (n_7718, n8640);
  and g16104 (n8641, n_7717, n_7718);
  not g16105 (n_7719, n8641);
  and g16106 (n8642, n8301, n_7719);
  not g16107 (n_7720, n8301);
  and g16108 (n8643, n_7720, n8641);
  not g16109 (n_7721, n8642);
  not g16110 (n_7722, n8643);
  and g16111 (n8644, n_7721, n_7722);
  and g16112 (n8645, n8204, n8317);
  not g16113 (n_7723, n8204);
  not g16114 (n_7724, n8317);
  and g16115 (n8646, n_7723, n_7724);
  not g16116 (n_7725, n8645);
  not g16117 (n_7726, n8646);
  and g16118 (n8647, n_7725, n_7726);
  not g16119 (n_7727, n8647);
  and g16120 (n8648, n8263, n_7727);
  not g16121 (n_7728, n8263);
  and g16122 (n8649, n_7728, n8647);
  not g16123 (n_7729, n8648);
  not g16124 (n_7730, n8649);
  and g16125 (n8650, n_7729, n_7730);
  and g16126 (n8651, n8644, n8650);
  not g16127 (n_7731, n8644);
  not g16128 (n_7732, n8650);
  and g16129 (n8652, n_7731, n_7732);
  not g16130 (n_7733, n8651);
  not g16131 (n_7734, n8652);
  and g16132 (n8653, n_7733, n_7734);
  not g16133 (n_7735, n8638);
  and g16134 (n8654, n_7735, n8653);
  not g16135 (n_7736, n8653);
  and g16136 (n8655, n8638, n_7736);
  not g16137 (n_7737, n8654);
  not g16138 (n_7738, n8655);
  and g16139 (n8656, n_7737, n_7738);
  not g16140 (n_7739, n8637);
  and g16141 (n8657, n_7739, n8656);
  not g16142 (n_7740, n8657);
  and g16143 (n8658, n_7739, n_7740);
  and g16144 (n8659, n8656, n_7740);
  not g16145 (n_7741, n8658);
  not g16146 (n_7742, n8659);
  and g16147 (n8660, n_7741, n_7742);
  not g16148 (n_7743, n8660);
  and g16149 (n8661, n8636, n_7743);
  not g16150 (n_7744, n8636);
  and g16151 (n8662, n_7744, n_7742);
  and g16152 (n8663, n_7741, n8662);
  not g16153 (n_7745, n8661);
  not g16154 (n_7746, n8663);
  and g16155 (n8664, n_7745, n_7746);
  not g16156 (n_7747, n8622);
  and g16157 (n8665, n_7747, n8664);
  not g16158 (n_7748, n8665);
  and g16159 (n8666, n_7747, n_7748);
  and g16160 (n8667, n8664, n_7748);
  not g16161 (n_7749, n8666);
  not g16162 (n_7750, n8667);
  and g16163 (n8668, n_7749, n_7750);
  not g16164 (n_7751, n8621);
  not g16165 (n_7752, n8668);
  and g16166 (n8669, n_7751, n_7752);
  and g16167 (n8670, n8621, n_7750);
  and g16168 (n8671, n_7749, n8670);
  not g16169 (n_7753, n8669);
  not g16170 (n_7754, n8671);
  and g16171 (n8672, n_7753, n_7754);
  and g16172 (n8673, n8432, n8672);
  not g16173 (n_7755, n8432);
  not g16174 (n_7756, n8672);
  and g16175 (n8674, n_7755, n_7756);
  not g16176 (n_7757, n8673);
  not g16177 (n_7758, n8674);
  and g16178 (n8675, n_7757, n_7758);
  not g16179 (n_7759, n8675);
  and g16180 (n8676, n8402, n_7759);
  not g16181 (n_7760, n8402);
  and g16182 (n8677, n_7760, n8675);
  not g16183 (n_7761, n8676);
  not g16184 (n_7762, n8677);
  and g16185 (n8678, n_7761, n_7762);
  and g16186 (n8679, n_7500, n_7504);
  not g16187 (n_7763, n8679);
  and g16188 (n8680, n_7501, n_7763);
  not g16189 (n_7764, n8678);
  and g16190 (n8681, n_7764, n8680);
  not g16191 (n_7765, n8680);
  and g16192 (n8682, n8678, n_7765);
  not g16193 (n_7766, n8681);
  not g16194 (n_7767, n8682);
  and g16195 (\asquared[61] , n_7766, n_7767);
  and g16196 (n8684, n_7535, n_7757);
  and g16197 (n8685, n_7748, n_7753);
  and g16198 (n8686, n_7613, n_7696);
  and g16199 (n8687, n_7710, n_7714);
  and g16200 (n8688, \a[7] , \a[54] );
  and g16201 (n8689, \a[8] , \a[53] );
  not g16202 (n_7768, n8688);
  not g16203 (n_7769, n8689);
  and g16204 (n8690, n_7768, n_7769);
  and g16205 (n8691, n380, n7699);
  not g16206 (n_7770, n8691);
  not g16209 (n_7771, n8690);
  not g16211 (n_7772, n8694);
  and g16212 (n8695, n_7770, n_7772);
  and g16213 (n8696, n_7771, n8695);
  and g16214 (n8697, \a[42] , n_7772);
  and g16215 (n8698, \a[19] , n8697);
  not g16216 (n_7773, n8696);
  not g16217 (n_7774, n8698);
  and g16218 (n8699, n_7773, n_7774);
  and g16219 (n8700, \a[44] , \a[52] );
  and g16220 (n8701, n1676, n8700);
  and g16221 (n8702, n6516, n8237);
  and g16222 (n8703, n1052, n5296);
  not g16223 (n_7775, n8702);
  not g16224 (n_7776, n8703);
  and g16225 (n8704, n_7775, n_7776);
  not g16226 (n_7777, n8701);
  not g16227 (n_7778, n8704);
  and g16228 (n8705, n_7777, n_7778);
  not g16229 (n_7779, n8705);
  and g16230 (n8706, \a[43] , n_7779);
  and g16231 (n8707, \a[18] , n8706);
  and g16232 (n8708, n_7777, n_7779);
  and g16233 (n8709, \a[9] , \a[52] );
  and g16234 (n8710, \a[17] , \a[44] );
  not g16235 (n_7780, n8709);
  not g16236 (n_7781, n8710);
  and g16237 (n8711, n_7780, n_7781);
  not g16238 (n_7782, n8711);
  and g16239 (n8712, n8708, n_7782);
  not g16240 (n_7783, n8707);
  not g16241 (n_7784, n8712);
  and g16242 (n8713, n_7783, n_7784);
  not g16243 (n_7785, n8699);
  not g16244 (n_7786, n8713);
  and g16245 (n8714, n_7785, n_7786);
  not g16246 (n_7787, n8714);
  and g16247 (n8715, n_7785, n_7787);
  and g16248 (n8716, n_7786, n_7787);
  not g16249 (n_7788, n8715);
  not g16250 (n_7789, n8716);
  and g16251 (n8717, n_7788, n_7789);
  and g16252 (n8718, n2331, n4150);
  and g16253 (n8719, n2800, n2972);
  and g16254 (n8720, n2227, n3319);
  not g16255 (n_7790, n8719);
  not g16256 (n_7791, n8720);
  and g16257 (n8721, n_7790, n_7791);
  not g16258 (n_7792, n8718);
  not g16259 (n_7793, n8721);
  and g16260 (n8722, n_7792, n_7793);
  not g16261 (n_7794, n8722);
  and g16262 (n8723, \a[35] , n_7794);
  and g16263 (n8724, \a[26] , n8723);
  and g16264 (n8725, n_7792, n_7794);
  and g16265 (n8726, \a[28] , \a[33] );
  not g16266 (n_7795, n3503);
  not g16267 (n_7796, n8726);
  and g16268 (n8727, n_7795, n_7796);
  not g16269 (n_7797, n8727);
  and g16270 (n8728, n8725, n_7797);
  not g16271 (n_7798, n8724);
  not g16272 (n_7799, n8728);
  and g16273 (n8729, n_7798, n_7799);
  not g16274 (n_7800, n8717);
  not g16275 (n_7801, n8729);
  and g16276 (n8730, n_7800, n_7801);
  not g16277 (n_7802, n8730);
  and g16278 (n8731, n_7800, n_7802);
  and g16279 (n8732, n_7801, n_7802);
  not g16280 (n_7803, n8731);
  not g16281 (n_7804, n8732);
  and g16282 (n8733, n_7803, n_7804);
  and g16283 (n8734, n_7733, n_7737);
  not g16284 (n_7805, n8733);
  not g16285 (n_7806, n8734);
  and g16286 (n8735, n_7805, n_7806);
  not g16287 (n_7807, n8735);
  and g16288 (n8736, n_7805, n_7807);
  and g16289 (n8737, n_7806, n_7807);
  not g16290 (n_7808, n8736);
  not g16291 (n_7809, n8737);
  and g16292 (n8738, n_7808, n_7809);
  not g16293 (n_7810, n8687);
  not g16294 (n_7811, n8738);
  and g16295 (n8739, n_7810, n_7811);
  not g16296 (n_7812, n8739);
  and g16297 (n8740, n_7810, n_7812);
  and g16298 (n8741, n_7811, n_7812);
  not g16299 (n_7813, n8740);
  not g16300 (n_7814, n8741);
  and g16301 (n8742, n_7813, n_7814);
  and g16302 (n8743, n_7579, n_7611);
  and g16303 (n8744, n_7726, n_7730);
  and g16304 (n8745, n_7702, n_7706);
  and g16305 (n8746, \a[3] , \a[58] );
  and g16306 (n8747, \a[4] , \a[57] );
  not g16307 (n_7815, n8746);
  not g16308 (n_7816, n8747);
  and g16309 (n8748, n_7815, n_7816);
  and g16310 (n8749, n209, n8436);
  not g16311 (n_7817, n8749);
  not g16314 (n_7818, n8748);
  not g16316 (n_7819, n8752);
  and g16317 (n8753, \a[38] , n_7819);
  and g16318 (n8754, \a[23] , n8753);
  and g16319 (n8755, n_7817, n_7819);
  and g16320 (n8756, n_7818, n8755);
  not g16321 (n_7820, n8754);
  not g16322 (n_7821, n8756);
  and g16323 (n8757, n_7820, n_7821);
  not g16324 (n_7822, n8745);
  not g16325 (n_7823, n8757);
  and g16326 (n8758, n_7822, n_7823);
  not g16327 (n_7824, n8758);
  and g16328 (n8759, n_7822, n_7824);
  and g16329 (n8760, n_7823, n_7824);
  not g16330 (n_7825, n8759);
  not g16331 (n_7826, n8760);
  and g16332 (n8761, n_7825, n_7826);
  not g16333 (n_7827, n8744);
  not g16334 (n_7828, n8761);
  and g16335 (n8762, n_7827, n_7828);
  not g16336 (n_7829, n8762);
  and g16337 (n8763, n_7827, n_7829);
  and g16338 (n8764, n_7828, n_7829);
  not g16339 (n_7830, n8763);
  not g16340 (n_7831, n8764);
  and g16341 (n8765, n_7830, n_7831);
  and g16342 (n8766, n_7591, n_7590);
  not g16343 (n_7832, n8766);
  and g16344 (n8767, n_7606, n_7832);
  and g16345 (n8768, n_7718, n_7722);
  and g16346 (n8769, \a[1] , \a[60] );
  and g16347 (n8770, \a[31] , n8769);
  not g16348 (n_7833, \a[31] );
  not g16349 (n_7834, n8769);
  and g16350 (n8771, n_7833, n_7834);
  not g16351 (n_7835, n8770);
  not g16352 (n_7836, n8771);
  and g16353 (n8772, n_7835, n_7836);
  and g16354 (n8773, n8535, n8772);
  not g16355 (n_7837, n8772);
  and g16356 (n8774, n_7620, n_7837);
  not g16357 (n_7838, n8773);
  not g16358 (n_7839, n8774);
  and g16359 (n8775, n_7838, n_7839);
  not g16360 (n_7840, n8584);
  and g16361 (n8776, n_7840, n8775);
  not g16362 (n_7841, n8775);
  and g16363 (n8777, n8584, n_7841);
  not g16364 (n_7842, n8776);
  not g16365 (n_7843, n8777);
  and g16366 (n8778, n_7842, n_7843);
  not g16367 (n_7844, n8768);
  and g16368 (n8779, n_7844, n8778);
  not g16369 (n_7845, n8778);
  and g16370 (n8780, n8768, n_7845);
  not g16371 (n_7846, n8779);
  not g16372 (n_7847, n8780);
  and g16373 (n8781, n_7846, n_7847);
  not g16374 (n_7848, n8767);
  and g16375 (n8782, n_7848, n8781);
  not g16376 (n_7849, n8781);
  and g16377 (n8783, n8767, n_7849);
  not g16378 (n_7850, n8782);
  not g16379 (n_7851, n8783);
  and g16380 (n8784, n_7850, n_7851);
  not g16381 (n_7852, n8765);
  and g16382 (n8785, n_7852, n8784);
  not g16383 (n_7853, n8785);
  and g16384 (n8786, n_7852, n_7853);
  and g16385 (n8787, n8784, n_7853);
  not g16386 (n_7854, n8786);
  not g16387 (n_7855, n8787);
  and g16388 (n8788, n_7854, n_7855);
  not g16389 (n_7856, n8743);
  not g16390 (n_7857, n8788);
  and g16391 (n8789, n_7856, n_7857);
  and g16392 (n8790, n8743, n_7855);
  and g16393 (n8791, n_7854, n8790);
  not g16394 (n_7858, n8789);
  not g16395 (n_7859, n8791);
  and g16396 (n8792, n_7858, n_7859);
  not g16397 (n_7860, n8742);
  and g16398 (n8793, n_7860, n8792);
  not g16399 (n_7861, n8793);
  and g16400 (n8794, n_7860, n_7861);
  and g16401 (n8795, n8792, n_7861);
  not g16402 (n_7862, n8794);
  not g16403 (n_7863, n8795);
  and g16404 (n8796, n_7862, n_7863);
  not g16405 (n_7864, n8686);
  not g16406 (n_7865, n8796);
  and g16407 (n8797, n_7864, n_7865);
  and g16408 (n8798, n8686, n_7863);
  and g16409 (n8799, n_7862, n8798);
  not g16410 (n_7866, n8797);
  not g16411 (n_7867, n8799);
  and g16412 (n8800, n_7866, n_7867);
  not g16413 (n_7868, n8685);
  and g16414 (n8801, n_7868, n8800);
  not g16415 (n_7869, n8801);
  and g16416 (n8802, n_7868, n_7869);
  and g16417 (n8803, n8800, n_7869);
  not g16418 (n_7870, n8802);
  not g16419 (n_7871, n8803);
  and g16420 (n8804, n_7870, n_7871);
  and g16421 (n8805, n_7690, n_7693);
  and g16422 (n8806, n8494, n8571);
  not g16423 (n_7872, n8494);
  not g16424 (n_7873, n8571);
  and g16425 (n8807, n_7872, n_7873);
  not g16426 (n_7874, n8806);
  not g16427 (n_7875, n8807);
  and g16428 (n8808, n_7874, n_7875);
  and g16429 (n8809, n_7617, n_7625);
  not g16430 (n_7876, n8808);
  and g16431 (n8810, n_7876, n8809);
  not g16432 (n_7877, n8809);
  and g16433 (n8811, n8808, n_7877);
  not g16434 (n_7878, n8810);
  not g16435 (n_7879, n8811);
  and g16436 (n8812, n_7878, n_7879);
  and g16437 (n8813, n_7669, n_7684);
  not g16438 (n_7880, n8812);
  and g16439 (n8814, n_7880, n8813);
  not g16440 (n_7881, n8813);
  and g16441 (n8815, n8812, n_7881);
  not g16442 (n_7882, n8814);
  not g16443 (n_7883, n8815);
  and g16444 (n8816, n_7882, n_7883);
  and g16445 (n8817, n_7640, n_7646);
  not g16446 (n_7884, n8816);
  and g16447 (n8818, n_7884, n8817);
  not g16448 (n_7885, n8817);
  and g16449 (n8819, n8816, n_7885);
  not g16450 (n_7886, n8818);
  not g16451 (n_7887, n8819);
  and g16452 (n8820, n_7886, n_7887);
  and g16453 (n8821, n_7558, n_7573);
  and g16454 (n8822, n8472, n8551);
  not g16455 (n_7888, n8472);
  not g16456 (n_7889, n8551);
  and g16457 (n8823, n_7888, n_7889);
  not g16458 (n_7890, n8822);
  not g16459 (n_7891, n8823);
  and g16460 (n8824, n_7890, n_7891);
  not g16461 (n_7892, n8824);
  and g16462 (n8825, n8458, n_7892);
  not g16463 (n_7893, n8458);
  and g16464 (n8826, n_7893, n8824);
  not g16465 (n_7894, n8825);
  not g16466 (n_7895, n8826);
  and g16467 (n8827, n_7894, n_7895);
  and g16468 (n8828, n8440, n8604);
  not g16469 (n_7896, n8440);
  not g16470 (n_7897, n8604);
  and g16471 (n8829, n_7896, n_7897);
  not g16472 (n_7898, n8828);
  not g16473 (n_7899, n8829);
  and g16474 (n8830, n_7898, n_7899);
  not g16475 (n_7900, n8830);
  and g16476 (n8831, n8515, n_7900);
  not g16477 (n_7901, n8515);
  and g16478 (n8832, n_7901, n8830);
  not g16479 (n_7902, n8831);
  not g16480 (n_7903, n8832);
  and g16481 (n8833, n_7902, n_7903);
  not g16482 (n_7904, n8827);
  not g16483 (n_7905, n8833);
  and g16484 (n8834, n_7904, n_7905);
  and g16485 (n8835, n8827, n8833);
  not g16486 (n_7906, n8834);
  not g16487 (n_7907, n8835);
  and g16488 (n8836, n_7906, n_7907);
  not g16489 (n_7908, n8821);
  and g16490 (n8837, n_7908, n8836);
  not g16491 (n_7909, n8836);
  and g16492 (n8838, n8821, n_7909);
  not g16493 (n_7910, n8837);
  not g16494 (n_7911, n8838);
  and g16495 (n8839, n_7910, n_7911);
  and g16496 (n8840, n8820, n8839);
  not g16497 (n_7912, n8820);
  not g16498 (n_7913, n8839);
  and g16499 (n8841, n_7912, n_7913);
  not g16500 (n_7914, n8805);
  not g16501 (n_7915, n8841);
  and g16502 (n8842, n_7914, n_7915);
  not g16503 (n_7916, n8840);
  and g16504 (n8843, n_7916, n8842);
  not g16505 (n_7917, n8843);
  and g16506 (n8844, n_7914, n_7917);
  and g16507 (n8845, n_7916, n_7917);
  and g16508 (n8846, n_7915, n8845);
  not g16509 (n_7918, n8844);
  not g16510 (n_7919, n8846);
  and g16511 (n8847, n_7918, n_7919);
  and g16512 (n8848, n_7526, n_7530);
  and g16513 (n8849, n8847, n8848);
  not g16514 (n_7920, n8847);
  not g16515 (n_7921, n8848);
  and g16516 (n8850, n_7920, n_7921);
  not g16517 (n_7922, n8849);
  not g16518 (n_7923, n8850);
  and g16519 (n8851, n_7922, n_7923);
  and g16520 (n8852, n_7740, n_7745);
  and g16521 (n8853, n_7519, n_7522);
  and g16522 (n8854, \a[46] , \a[51] );
  and g16523 (n8855, n685, n8854);
  and g16524 (n8856, n891, n5560);
  and g16525 (n8857, \a[10] , \a[51] );
  and g16526 (n8858, n5850, n8857);
  not g16527 (n_7924, n8856);
  not g16528 (n_7925, n8858);
  and g16529 (n8859, n_7924, n_7925);
  not g16530 (n_7926, n8855);
  not g16531 (n_7927, n8859);
  and g16532 (n8860, n_7926, n_7927);
  not g16533 (n_7928, n8860);
  and g16534 (n8861, n_7926, n_7928);
  and g16535 (n8862, \a[15] , \a[46] );
  not g16536 (n_7929, n8857);
  not g16537 (n_7930, n8862);
  and g16538 (n8863, n_7929, n_7930);
  not g16539 (n_7931, n8863);
  and g16540 (n8864, n8861, n_7931);
  and g16541 (n8865, n5850, n_7928);
  not g16542 (n_7932, n8864);
  not g16543 (n_7933, n8865);
  and g16544 (n8866, n_7932, n_7933);
  and g16545 (n8867, n606, n6254);
  and g16546 (n8868, \a[14] , \a[50] );
  and g16547 (n8869, n8060, n8868);
  and g16548 (n8870, n602, n6325);
  not g16549 (n_7934, n8869);
  not g16550 (n_7935, n8870);
  and g16551 (n8871, n_7934, n_7935);
  not g16552 (n_7936, n8867);
  not g16553 (n_7937, n8871);
  and g16554 (n8872, n_7936, n_7937);
  not g16555 (n_7938, n8872);
  and g16556 (n8873, \a[50] , n_7938);
  and g16557 (n8874, \a[11] , n8873);
  and g16558 (n8875, n_7936, n_7938);
  and g16559 (n8876, \a[12] , \a[49] );
  not g16560 (n_7939, n7403);
  not g16561 (n_7940, n8876);
  and g16562 (n8877, n_7939, n_7940);
  not g16563 (n_7941, n8877);
  and g16564 (n8878, n8875, n_7941);
  not g16565 (n_7942, n8874);
  not g16566 (n_7943, n8878);
  and g16567 (n8879, n_7942, n_7943);
  not g16568 (n_7944, n8866);
  not g16569 (n_7945, n8879);
  and g16570 (n8880, n_7944, n_7945);
  not g16571 (n_7946, n8880);
  and g16572 (n8881, n_7944, n_7946);
  and g16573 (n8882, n_7945, n_7946);
  not g16574 (n_7947, n8881);
  not g16575 (n_7948, n8882);
  and g16576 (n8883, n_7947, n_7948);
  and g16577 (n8884, \a[29] , \a[32] );
  not g16578 (n_7949, n2865);
  not g16579 (n_7950, n8884);
  and g16580 (n8885, n_7949, n_7950);
  and g16581 (n8886, n2617, n3812);
  not g16582 (n_7951, n8886);
  not g16585 (n_7952, n8885);
  not g16587 (n_7953, n8889);
  and g16588 (n8890, \a[48] , n_7953);
  and g16589 (n8891, \a[13] , n8890);
  and g16590 (n8892, n_7951, n_7953);
  and g16591 (n8893, n_7952, n8892);
  not g16592 (n_7954, n8891);
  not g16593 (n_7955, n8893);
  and g16594 (n8894, n_7954, n_7955);
  not g16595 (n_7956, n8883);
  not g16596 (n_7957, n8894);
  and g16597 (n8895, n_7956, n_7957);
  not g16598 (n_7958, n8895);
  and g16599 (n8896, n_7956, n_7958);
  and g16600 (n8897, n_7957, n_7958);
  not g16601 (n_7959, n8896);
  not g16602 (n_7960, n8897);
  and g16603 (n8898, n_7959, n_7960);
  and g16604 (n8899, n_7510, n_7515);
  and g16605 (n8900, n8898, n8899);
  not g16606 (n_7961, n8898);
  not g16607 (n_7962, n8899);
  and g16608 (n8901, n_7961, n_7962);
  not g16609 (n_7963, n8900);
  not g16610 (n_7964, n8901);
  and g16611 (n8902, n_7963, n_7964);
  and g16612 (n8903, \a[5] , \a[59] );
  and g16613 (n8904, n7953, n8903);
  and g16614 (n8905, \a[59] , \a[61] );
  and g16615 (n8906, n196, n8905);
  and g16616 (n8907, \a[5] , \a[61] );
  and g16617 (n8908, n7423, n8907);
  not g16618 (n_7966, n8906);
  not g16619 (n_7967, n8908);
  and g16620 (n8909, n_7966, n_7967);
  not g16621 (n_7968, n8904);
  not g16622 (n_7969, n8909);
  and g16623 (n8910, n_7968, n_7969);
  not g16624 (n_7970, n8910);
  and g16625 (n8911, n_7968, n_7970);
  and g16626 (n8912, \a[2] , \a[59] );
  and g16627 (n8913, \a[5] , \a[56] );
  not g16628 (n_7971, n8912);
  not g16629 (n_7972, n8913);
  and g16630 (n8914, n_7971, n_7972);
  not g16631 (n_7973, n8914);
  and g16632 (n8915, n8911, n_7973);
  and g16633 (n8916, \a[61] , n_7970);
  and g16634 (n8917, \a[0] , n8916);
  not g16635 (n_7974, n8915);
  not g16636 (n_7975, n8917);
  and g16637 (n8918, n_7974, n_7975);
  and g16638 (n8919, \a[20] , \a[41] );
  and g16639 (n8920, \a[21] , \a[40] );
  not g16640 (n_7976, n8919);
  not g16641 (n_7977, n8920);
  and g16642 (n8921, n_7976, n_7977);
  and g16643 (n8922, n1494, n5413);
  not g16644 (n_7978, n8922);
  not g16647 (n_7979, n8921);
  not g16649 (n_7980, n8925);
  and g16650 (n8926, \a[55] , n_7980);
  and g16651 (n8927, \a[6] , n8926);
  and g16652 (n8928, n_7978, n_7980);
  and g16653 (n8929, n_7979, n8928);
  not g16654 (n_7981, n8927);
  not g16655 (n_7982, n8929);
  and g16656 (n8930, n_7981, n_7982);
  not g16657 (n_7983, n8918);
  not g16658 (n_7984, n8930);
  and g16659 (n8931, n_7983, n_7984);
  not g16660 (n_7985, n8931);
  and g16661 (n8932, n_7983, n_7985);
  and g16662 (n8933, n_7984, n_7985);
  not g16663 (n_7986, n8932);
  not g16664 (n_7987, n8933);
  and g16665 (n8934, n_7986, n_7987);
  and g16666 (n8935, n1904, n3687);
  and g16667 (n8936, \a[36] , \a[39] );
  and g16668 (n8937, n5327, n8936);
  and g16669 (n8938, n2115, n5430);
  not g16670 (n_7988, n8937);
  not g16671 (n_7989, n8938);
  and g16672 (n8939, n_7988, n_7989);
  not g16673 (n_7990, n8935);
  not g16674 (n_7991, n8939);
  and g16675 (n8940, n_7990, n_7991);
  not g16676 (n_7992, n8940);
  and g16677 (n8941, \a[39] , n_7992);
  and g16678 (n8942, \a[22] , n8941);
  and g16679 (n8943, \a[24] , \a[37] );
  and g16680 (n8944, \a[25] , \a[36] );
  not g16681 (n_7993, n8943);
  not g16682 (n_7994, n8944);
  and g16683 (n8945, n_7993, n_7994);
  and g16684 (n8946, n_7990, n_7992);
  not g16685 (n_7995, n8945);
  and g16686 (n8947, n_7995, n8946);
  not g16687 (n_7996, n8942);
  not g16688 (n_7997, n8947);
  and g16689 (n8948, n_7996, n_7997);
  not g16690 (n_7998, n8934);
  not g16691 (n_7999, n8948);
  and g16692 (n8949, n_7998, n_7999);
  not g16693 (n_8000, n8949);
  and g16694 (n8950, n_7998, n_8000);
  and g16695 (n8951, n_7999, n_8000);
  not g16696 (n_8001, n8950);
  not g16697 (n_8002, n8951);
  and g16698 (n8952, n_8001, n_8002);
  not g16699 (n_8003, n8902);
  and g16700 (n8953, n_8003, n8952);
  not g16701 (n_8004, n8952);
  and g16702 (n8954, n8902, n_8004);
  not g16703 (n_8005, n8953);
  not g16704 (n_8006, n8954);
  and g16705 (n8955, n_8005, n_8006);
  not g16706 (n_8007, n8853);
  and g16707 (n8956, n_8007, n8955);
  not g16708 (n_8008, n8955);
  and g16709 (n8957, n8853, n_8008);
  not g16710 (n_8009, n8956);
  not g16711 (n_8010, n8957);
  and g16712 (n8958, n_8009, n_8010);
  not g16713 (n_8011, n8852);
  and g16714 (n8959, n_8011, n8958);
  not g16715 (n_8012, n8958);
  and g16716 (n8960, n8852, n_8012);
  not g16717 (n_8013, n8959);
  not g16718 (n_8014, n8960);
  and g16719 (n8961, n_8013, n_8014);
  and g16720 (n8962, n8851, n8961);
  not g16721 (n_8015, n8851);
  not g16722 (n_8016, n8961);
  and g16723 (n8963, n_8015, n_8016);
  not g16724 (n_8017, n8962);
  not g16725 (n_8018, n8963);
  and g16726 (n8964, n_8017, n_8018);
  not g16727 (n_8019, n8804);
  and g16728 (n8965, n_8019, n8964);
  not g16729 (n_8020, n8964);
  and g16730 (n8966, n_7871, n_8020);
  and g16731 (n8967, n_7870, n8966);
  not g16732 (n_8021, n8965);
  not g16733 (n_8022, n8967);
  and g16734 (n8968, n_8021, n_8022);
  not g16735 (n_8023, n8684);
  and g16736 (n8969, n_8023, n8968);
  not g16737 (n_8024, n8968);
  and g16738 (n8970, n8684, n_8024);
  not g16739 (n_8025, n8969);
  not g16740 (n_8026, n8970);
  and g16741 (n8971, n_8025, n_8026);
  and g16742 (n8972, n_7761, n_7765);
  not g16743 (n_8027, n8972);
  and g16744 (n8973, n_7762, n_8027);
  not g16745 (n_8028, n8971);
  and g16746 (n8974, n_8028, n8973);
  not g16747 (n_8029, n8973);
  and g16748 (n8975, n8971, n_8029);
  not g16749 (n_8030, n8974);
  not g16750 (n_8031, n8975);
  and g16751 (\asquared[62] , n_8030, n_8031);
  and g16752 (n8977, n_8026, n_8029);
  not g16753 (n_8032, n8977);
  and g16754 (n8978, n_8025, n_8032);
  and g16755 (n8979, n_7869, n_8021);
  and g16756 (n8980, n_7861, n_7866);
  and g16757 (n8981, n8708, n8861);
  not g16758 (n_8033, n8708);
  not g16759 (n_8034, n8861);
  and g16760 (n8982, n_8033, n_8034);
  not g16761 (n_8035, n8981);
  not g16762 (n_8036, n8982);
  and g16763 (n8983, n_8035, n_8036);
  and g16764 (n8984, n226, n8436);
  and g16765 (n8985, \a[57] , \a[59] );
  and g16766 (n8986, n300, n8985);
  and g16767 (n8987, \a[58] , \a[59] );
  and g16768 (n8988, n209, n8987);
  not g16769 (n_8037, n8986);
  not g16770 (n_8038, n8988);
  and g16771 (n8989, n_8037, n_8038);
  not g16772 (n_8039, n8984);
  not g16773 (n_8040, n8989);
  and g16774 (n8990, n_8039, n_8040);
  not g16775 (n_8041, n8990);
  and g16776 (n8991, \a[59] , n_8041);
  and g16777 (n8992, \a[3] , n8991);
  and g16778 (n8993, n_8039, n_8041);
  and g16779 (n8994, \a[4] , \a[58] );
  and g16780 (n8995, \a[5] , \a[57] );
  not g16781 (n_8042, n8994);
  not g16782 (n_8043, n8995);
  and g16783 (n8996, n_8042, n_8043);
  not g16784 (n_8044, n8996);
  and g16785 (n8997, n8993, n_8044);
  not g16786 (n_8045, n8992);
  not g16787 (n_8046, n8997);
  and g16788 (n8998, n_8045, n_8046);
  not g16789 (n_8047, n8998);
  and g16790 (n8999, n8983, n_8047);
  not g16791 (n_8048, n8999);
  and g16792 (n9000, n8983, n_8048);
  and g16793 (n9001, n_8047, n_8048);
  not g16794 (n_8049, n9000);
  not g16795 (n_8050, n9001);
  and g16796 (n9002, n_8049, n_8050);
  and g16797 (n9003, n_7787, n_7802);
  and g16798 (n9004, n9002, n9003);
  not g16799 (n_8051, n9002);
  not g16800 (n_8052, n9003);
  and g16801 (n9005, n_8051, n_8052);
  not g16802 (n_8053, n9004);
  not g16803 (n_8054, n9005);
  and g16804 (n9006, n_8053, n_8054);
  and g16805 (n9007, n_7824, n_7829);
  not g16806 (n_8055, n9006);
  and g16807 (n9008, n_8055, n9007);
  not g16808 (n_8056, n9007);
  and g16809 (n9009, n9006, n_8056);
  not g16810 (n_8057, n9008);
  not g16811 (n_8058, n9009);
  and g16812 (n9010, n_8057, n_8058);
  and g16813 (n9011, n_7875, n_7879);
  and g16814 (n9012, n_7838, n_7842);
  and g16815 (n9013, n9011, n9012);
  not g16816 (n_8059, n9011);
  not g16817 (n_8060, n9012);
  and g16818 (n9014, n_8059, n_8060);
  not g16819 (n_8061, n9013);
  not g16820 (n_8062, n9014);
  and g16821 (n9015, n_8061, n_8062);
  and g16822 (n9016, n_7891, n_7895);
  not g16823 (n_8063, n9015);
  and g16824 (n9017, n_8063, n9016);
  not g16825 (n_8064, n9016);
  and g16826 (n9018, n9015, n_8064);
  not g16827 (n_8065, n9017);
  not g16828 (n_8066, n9018);
  and g16829 (n9019, n_8065, n_8066);
  and g16830 (n9020, n_7964, n_8006);
  not g16831 (n_8067, n9020);
  and g16832 (n9021, n9019, n_8067);
  not g16833 (n_8068, n9021);
  and g16834 (n9022, n9019, n_8068);
  and g16835 (n9023, n_8067, n_8068);
  not g16836 (n_8069, n9022);
  not g16837 (n_8070, n9023);
  and g16838 (n9024, n_8069, n_8070);
  not g16839 (n_8071, n9024);
  and g16840 (n9025, n9010, n_8071);
  not g16841 (n_8072, n9010);
  and g16842 (n9026, n_8072, n_8070);
  and g16843 (n9027, n_8069, n9026);
  not g16844 (n_8073, n9025);
  not g16845 (n_8074, n9027);
  and g16846 (n9028, n_8073, n_8074);
  not g16847 (n_8075, n8980);
  and g16848 (n9029, n_8075, n9028);
  not g16849 (n_8076, n9028);
  and g16850 (n9030, n8980, n_8076);
  not g16851 (n_8077, n9029);
  not g16852 (n_8078, n9030);
  and g16853 (n9031, n_8077, n_8078);
  and g16854 (n9032, n_7853, n_7858);
  and g16855 (n9033, \a[8] , \a[54] );
  and g16856 (n9034, \a[18] , \a[44] );
  not g16857 (n_8079, n9033);
  not g16858 (n_8080, n9034);
  and g16859 (n9035, n_8079, n_8080);
  and g16860 (n9036, \a[18] , \a[54] );
  and g16861 (n9037, n6469, n9036);
  and g16862 (n9038, n1149, n5296);
  and g16863 (n9039, \a[19] , \a[54] );
  and g16864 (n9040, n6173, n9039);
  not g16865 (n_8081, n9038);
  not g16866 (n_8082, n9040);
  and g16867 (n9041, n_8081, n_8082);
  not g16868 (n_8083, n9037);
  not g16869 (n_8084, n9041);
  and g16870 (n9042, n_8083, n_8084);
  not g16871 (n_8085, n9042);
  and g16872 (n9043, n_8083, n_8085);
  not g16873 (n_8086, n9035);
  and g16874 (n9044, n_8086, n9043);
  and g16875 (n9045, \a[43] , n_8085);
  and g16876 (n9046, \a[19] , n9045);
  not g16877 (n_8087, n9044);
  not g16878 (n_8088, n9046);
  and g16879 (n9047, n_8087, n_8088);
  and g16880 (n9048, n2334, n4150);
  and g16881 (n9049, n2041, n2972);
  and g16882 (n9050, n2331, n3319);
  not g16883 (n_8089, n9049);
  not g16884 (n_8090, n9050);
  and g16885 (n9051, n_8089, n_8090);
  not g16886 (n_8091, n9048);
  not g16887 (n_8092, n9051);
  and g16888 (n9052, n_8091, n_8092);
  not g16889 (n_8093, n9052);
  and g16890 (n9053, \a[35] , n_8093);
  and g16891 (n9054, \a[27] , n9053);
  and g16892 (n9055, n_8091, n_8093);
  and g16893 (n9056, \a[28] , \a[34] );
  and g16894 (n9057, \a[29] , \a[33] );
  not g16895 (n_8094, n9056);
  not g16896 (n_8095, n9057);
  and g16897 (n9058, n_8094, n_8095);
  not g16898 (n_8096, n9058);
  and g16899 (n9059, n9055, n_8096);
  not g16900 (n_8097, n9054);
  not g16901 (n_8098, n9059);
  and g16902 (n9060, n_8097, n_8098);
  not g16903 (n_8099, n9047);
  not g16904 (n_8100, n9060);
  and g16905 (n9061, n_8099, n_8100);
  not g16906 (n_8101, n9061);
  and g16907 (n9062, n_8099, n_8101);
  and g16908 (n9063, n_8100, n_8101);
  not g16909 (n_8102, n9062);
  not g16910 (n_8103, n9063);
  and g16911 (n9064, n_8102, n_8103);
  and g16912 (n9065, n1666, n5083);
  and g16913 (n9066, n2115, n3803);
  and g16914 (n9067, n1919, n4171);
  not g16915 (n_8104, n9066);
  not g16916 (n_8105, n9067);
  and g16917 (n9068, n_8104, n_8105);
  not g16918 (n_8106, n9065);
  not g16919 (n_8107, n9068);
  and g16920 (n9069, n_8106, n_8107);
  not g16921 (n_8108, n9069);
  and g16922 (n9070, \a[40] , n_8108);
  and g16923 (n9071, \a[22] , n9070);
  and g16924 (n9072, n_8106, n_8108);
  and g16925 (n9073, \a[23] , \a[39] );
  and g16926 (n9074, \a[24] , \a[38] );
  not g16927 (n_8109, n9073);
  not g16928 (n_8110, n9074);
  and g16929 (n9075, n_8109, n_8110);
  not g16930 (n_8111, n9075);
  and g16931 (n9076, n9072, n_8111);
  not g16932 (n_8112, n9071);
  not g16933 (n_8113, n9076);
  and g16934 (n9077, n_8112, n_8113);
  not g16935 (n_8114, n9064);
  not g16936 (n_8115, n9077);
  and g16937 (n9078, n_8114, n_8115);
  not g16938 (n_8116, n9078);
  and g16939 (n9079, n_8114, n_8116);
  and g16940 (n9080, n_8115, n_8116);
  not g16941 (n_8117, n9079);
  not g16942 (n_8118, n9080);
  and g16943 (n9081, n_8117, n_8118);
  and g16944 (n9082, \a[0] , \a[62] );
  and g16945 (n9083, \a[2] , \a[60] );
  not g16946 (n_8120, n9082);
  not g16947 (n_8121, n9083);
  and g16948 (n9084, n_8120, n_8121);
  and g16949 (n9085, \a[60] , \a[62] );
  and g16950 (n9086, n196, n9085);
  not g16951 (n_8122, n9084);
  not g16952 (n_8123, n9086);
  and g16953 (n9087, n_8122, n_8123);
  and g16954 (n9088, n8770, n9087);
  not g16955 (n_8124, n9088);
  and g16956 (n9089, n_8123, n_8124);
  and g16957 (n9090, n_8122, n9089);
  and g16958 (n9091, n8770, n_8124);
  not g16959 (n_8125, n9090);
  not g16960 (n_8126, n9091);
  and g16961 (n9092, n_8125, n_8126);
  and g16962 (n9093, \a[21] , \a[41] );
  and g16963 (n9094, \a[25] , \a[37] );
  and g16964 (n9095, \a[26] , \a[36] );
  not g16965 (n_8127, n9094);
  not g16966 (n_8128, n9095);
  and g16967 (n9096, n_8127, n_8128);
  and g16968 (n9097, n2463, n3687);
  not g16969 (n_8129, n9097);
  and g16970 (n9098, n9093, n_8129);
  not g16971 (n_8130, n9096);
  and g16972 (n9099, n_8130, n9098);
  not g16973 (n_8131, n9099);
  and g16974 (n9100, n9093, n_8131);
  and g16975 (n9101, n_8129, n_8131);
  and g16976 (n9102, n_8130, n9101);
  not g16977 (n_8132, n9100);
  not g16978 (n_8133, n9102);
  and g16979 (n9103, n_8132, n_8133);
  not g16980 (n_8134, n9092);
  not g16981 (n_8135, n9103);
  and g16982 (n9104, n_8134, n_8135);
  not g16983 (n_8136, n9104);
  and g16984 (n9105, n_8134, n_8136);
  and g16985 (n9106, n_8135, n_8136);
  not g16986 (n_8137, n9105);
  not g16987 (n_8138, n9106);
  and g16988 (n9107, n_8137, n_8138);
  and g16989 (n9108, \a[45] , \a[52] );
  and g16990 (n9109, n1858, n9108);
  and g16991 (n9110, n484, n7433);
  and g16992 (n9111, \a[17] , \a[53] );
  and g16993 (n9112, n6997, n9111);
  not g16994 (n_8139, n9110);
  not g16995 (n_8140, n9112);
  and g16996 (n9113, n_8139, n_8140);
  not g16997 (n_8141, n9109);
  not g16998 (n_8142, n9113);
  and g16999 (n9114, n_8141, n_8142);
  not g17000 (n_8143, n9114);
  and g17001 (n9115, \a[53] , n_8143);
  and g17002 (n9116, \a[9] , n9115);
  and g17003 (n9117, n_8141, n_8143);
  and g17004 (n9118, \a[10] , \a[52] );
  and g17005 (n9119, \a[17] , \a[45] );
  not g17006 (n_8144, n9118);
  not g17007 (n_8145, n9119);
  and g17008 (n9120, n_8144, n_8145);
  not g17009 (n_8146, n9120);
  and g17010 (n9121, n9117, n_8146);
  not g17011 (n_8147, n9116);
  not g17012 (n_8148, n9121);
  and g17013 (n9122, n_8147, n_8148);
  not g17014 (n_8149, n9107);
  not g17015 (n_8150, n9122);
  and g17016 (n9123, n_8149, n_8150);
  not g17017 (n_8151, n9123);
  and g17018 (n9124, n_8149, n_8151);
  and g17019 (n9125, n_8150, n_8151);
  not g17020 (n_8152, n9124);
  not g17021 (n_8153, n9125);
  and g17022 (n9126, n_8152, n_8153);
  and g17023 (n9127, \a[47] , \a[51] );
  and g17024 (n9128, n816, n9127);
  and g17025 (n9129, n1843, n8854);
  and g17026 (n9130, n891, n5666);
  not g17027 (n_8154, n9129);
  not g17028 (n_8155, n9130);
  and g17029 (n9131, n_8154, n_8155);
  not g17030 (n_8156, n9128);
  not g17031 (n_8157, n9131);
  and g17032 (n9132, n_8156, n_8157);
  not g17033 (n_8158, n9132);
  and g17034 (n9133, n_8156, n_8158);
  and g17035 (n9134, \a[11] , \a[51] );
  and g17036 (n9135, \a[15] , \a[47] );
  not g17037 (n_8159, n9134);
  not g17038 (n_8160, n9135);
  and g17039 (n9136, n_8159, n_8160);
  not g17040 (n_8161, n9136);
  and g17041 (n9137, n9133, n_8161);
  and g17042 (n9138, \a[46] , n_8158);
  and g17043 (n9139, \a[16] , n9138);
  not g17044 (n_8162, n9137);
  not g17045 (n_8163, n9139);
  and g17046 (n9140, n_8162, n_8163);
  and g17047 (n9141, n745, n6256);
  and g17048 (n9142, n606, n5888);
  and g17049 (n9143, n748, n6325);
  not g17050 (n_8164, n9142);
  not g17051 (n_8165, n9143);
  and g17052 (n9144, n_8164, n_8165);
  not g17053 (n_8166, n9141);
  not g17054 (n_8167, n9144);
  and g17055 (n9145, n_8166, n_8167);
  not g17056 (n_8168, n9145);
  and g17057 (n9146, \a[50] , n_8168);
  and g17058 (n9147, \a[12] , n9146);
  and g17059 (n9148, \a[13] , \a[49] );
  and g17060 (n9149, \a[14] , \a[48] );
  not g17061 (n_8169, n9148);
  not g17062 (n_8170, n9149);
  and g17063 (n9150, n_8169, n_8170);
  and g17064 (n9151, n_8166, n_8168);
  not g17065 (n_8171, n9150);
  and g17066 (n9152, n_8171, n9151);
  not g17067 (n_8172, n9147);
  not g17068 (n_8173, n9152);
  and g17069 (n9153, n_8172, n_8173);
  not g17070 (n_8174, n9140);
  not g17071 (n_8175, n9153);
  and g17072 (n9154, n_8174, n_8175);
  not g17073 (n_8176, n9154);
  and g17074 (n9155, n_8174, n_8176);
  and g17075 (n9156, n_8175, n_8176);
  not g17076 (n_8177, n9155);
  not g17077 (n_8178, n9156);
  and g17078 (n9157, n_8177, n_8178);
  and g17079 (n9158, \a[6] , \a[56] );
  and g17080 (n9159, \a[7] , \a[55] );
  not g17081 (n_8179, n9158);
  not g17082 (n_8180, n9159);
  and g17083 (n9160, n_8179, n_8180);
  and g17084 (n9161, \a[55] , \a[56] );
  and g17085 (n9162, n335, n9161);
  not g17086 (n_8181, n9162);
  not g17089 (n_8182, n9160);
  not g17091 (n_8183, n9165);
  and g17092 (n9166, \a[42] , n_8183);
  and g17093 (n9167, \a[20] , n9166);
  and g17094 (n9168, n_8181, n_8183);
  and g17095 (n9169, n_8182, n9168);
  not g17096 (n_8184, n9167);
  not g17097 (n_8185, n9169);
  and g17098 (n9170, n_8184, n_8185);
  not g17099 (n_8186, n9157);
  not g17100 (n_8187, n9170);
  and g17101 (n9171, n_8186, n_8187);
  not g17102 (n_8188, n9171);
  and g17103 (n9172, n_8186, n_8188);
  and g17104 (n9173, n_8187, n_8188);
  not g17105 (n_8189, n9172);
  not g17106 (n_8190, n9173);
  and g17107 (n9174, n_8189, n_8190);
  not g17108 (n_8191, n9126);
  and g17109 (n9175, n_8191, n9174);
  not g17110 (n_8192, n9174);
  and g17111 (n9176, n9126, n_8192);
  not g17112 (n_8193, n9175);
  not g17113 (n_8194, n9176);
  and g17114 (n9177, n_8193, n_8194);
  not g17115 (n_8195, n9081);
  not g17116 (n_8196, n9177);
  and g17117 (n9178, n_8195, n_8196);
  and g17118 (n9179, n9081, n9177);
  not g17119 (n_8197, n9178);
  not g17120 (n_8198, n9179);
  and g17121 (n9180, n_8197, n_8198);
  not g17122 (n_8199, n9032);
  and g17123 (n9181, n_8199, n9180);
  not g17124 (n_8200, n9181);
  and g17125 (n9182, n_8199, n_8200);
  and g17126 (n9183, n9180, n_8200);
  not g17127 (n_8201, n9182);
  not g17128 (n_8202, n9183);
  and g17129 (n9184, n_8201, n_8202);
  not g17130 (n_8203, n8845);
  not g17131 (n_8204, n9184);
  and g17132 (n9185, n_8203, n_8204);
  not g17133 (n_8205, n9185);
  and g17134 (n9186, n_8203, n_8205);
  and g17135 (n9187, n_8204, n_8205);
  not g17136 (n_8206, n9186);
  not g17137 (n_8207, n9187);
  and g17138 (n9188, n_8206, n_8207);
  not g17139 (n_8208, n9031);
  and g17140 (n9189, n_8208, n9188);
  not g17141 (n_8209, n9188);
  and g17142 (n9190, n9031, n_8209);
  not g17143 (n_8210, n9189);
  not g17144 (n_8211, n9190);
  and g17145 (n9191, n_8210, n_8211);
  and g17146 (n9192, n_7923, n_8017);
  and g17147 (n9193, n_7899, n_7903);
  and g17148 (n9194, n_7985, n_8000);
  and g17149 (n9195, n9193, n9194);
  not g17150 (n_8212, n9193);
  not g17151 (n_8213, n9194);
  and g17152 (n9196, n_8212, n_8213);
  not g17153 (n_8214, n9195);
  not g17154 (n_8215, n9196);
  and g17155 (n9197, n_8214, n_8215);
  and g17156 (n9198, n_7946, n_7958);
  not g17157 (n_8216, n9197);
  and g17158 (n9199, n_8216, n9198);
  not g17159 (n_8217, n9198);
  and g17160 (n9200, n9197, n_8217);
  not g17161 (n_8218, n9199);
  not g17162 (n_8219, n9200);
  and g17163 (n9201, n_8218, n_8219);
  and g17164 (n9202, n8911, n8928);
  not g17165 (n_8220, n8911);
  not g17166 (n_8221, n8928);
  and g17167 (n9203, n_8220, n_8221);
  not g17168 (n_8222, n9202);
  not g17169 (n_8223, n9203);
  and g17170 (n9204, n_8222, n_8223);
  not g17171 (n_8224, n9204);
  and g17172 (n9205, n8695, n_8224);
  not g17173 (n_8225, n8695);
  and g17174 (n9206, n_8225, n9204);
  not g17175 (n_8226, n9205);
  not g17176 (n_8227, n9206);
  and g17177 (n9207, n_8226, n_8227);
  and g17178 (n9208, n8725, n8755);
  not g17179 (n_8228, n8725);
  not g17180 (n_8229, n8755);
  and g17181 (n9209, n_8228, n_8229);
  not g17182 (n_8230, n9208);
  not g17183 (n_8231, n9209);
  and g17184 (n9210, n_8230, n_8231);
  not g17185 (n_8232, n9210);
  and g17186 (n9211, n8946, n_8232);
  not g17187 (n_8233, n8946);
  and g17188 (n9212, n_8233, n9210);
  not g17189 (n_8234, n9211);
  not g17190 (n_8235, n9212);
  and g17191 (n9213, n_8234, n_8235);
  and g17192 (n9214, \a[1] , \a[61] );
  and g17193 (n9215, n2488, n9214);
  not g17194 (n_8236, n2488);
  not g17195 (n_8237, n9214);
  and g17196 (n9216, n_8236, n_8237);
  not g17197 (n_8238, n9215);
  not g17198 (n_8239, n9216);
  and g17199 (n9217, n_8238, n_8239);
  not g17200 (n_8240, n9217);
  and g17201 (n9218, n8892, n_8240);
  not g17202 (n_8241, n8892);
  and g17203 (n9219, n_8241, n9217);
  not g17204 (n_8242, n9218);
  not g17205 (n_8243, n9219);
  and g17206 (n9220, n_8242, n_8243);
  not g17207 (n_8244, n8875);
  and g17208 (n9221, n_8244, n9220);
  not g17209 (n_8245, n9220);
  and g17210 (n9222, n8875, n_8245);
  not g17211 (n_8246, n9221);
  not g17212 (n_8247, n9222);
  and g17213 (n9223, n_8246, n_8247);
  and g17214 (n9224, n9213, n9223);
  not g17215 (n_8248, n9224);
  and g17216 (n9225, n9213, n_8248);
  and g17217 (n9226, n9223, n_8248);
  not g17218 (n_8249, n9225);
  not g17219 (n_8250, n9226);
  and g17220 (n9227, n_8249, n_8250);
  not g17221 (n_8251, n9227);
  and g17222 (n9228, n9207, n_8251);
  not g17223 (n_8252, n9228);
  and g17224 (n9229, n9207, n_8252);
  and g17225 (n9230, n_8251, n_8252);
  not g17226 (n_8253, n9229);
  not g17227 (n_8254, n9230);
  and g17228 (n9231, n_8253, n_8254);
  not g17229 (n_8255, n9231);
  and g17230 (n9232, n9201, n_8255);
  not g17231 (n_8256, n9232);
  and g17232 (n9233, n9201, n_8256);
  and g17233 (n9234, n_8255, n_8256);
  not g17234 (n_8257, n9233);
  not g17235 (n_8258, n9234);
  and g17236 (n9235, n_8257, n_8258);
  and g17237 (n9236, n_7807, n_7812);
  and g17238 (n9237, n9235, n9236);
  not g17239 (n_8259, n9235);
  not g17240 (n_8260, n9236);
  and g17241 (n9238, n_8259, n_8260);
  not g17242 (n_8261, n9237);
  not g17243 (n_8262, n9238);
  and g17244 (n9239, n_8261, n_8262);
  and g17245 (n9240, n_7907, n_7910);
  and g17246 (n9241, n_7846, n_7850);
  and g17247 (n9242, n9240, n9241);
  not g17248 (n_8263, n9240);
  not g17249 (n_8264, n9241);
  and g17250 (n9243, n_8263, n_8264);
  not g17251 (n_8265, n9242);
  not g17252 (n_8266, n9243);
  and g17253 (n9244, n_8265, n_8266);
  and g17254 (n9245, n_7883, n_7887);
  not g17255 (n_8267, n9244);
  and g17256 (n9246, n_8267, n9245);
  not g17257 (n_8268, n9245);
  and g17258 (n9247, n9244, n_8268);
  not g17259 (n_8269, n9246);
  not g17260 (n_8270, n9247);
  and g17261 (n9248, n_8269, n_8270);
  and g17262 (n9249, n_8009, n_8013);
  not g17263 (n_8271, n9248);
  and g17264 (n9250, n_8271, n9249);
  not g17265 (n_8272, n9249);
  and g17266 (n9251, n9248, n_8272);
  not g17267 (n_8273, n9250);
  not g17268 (n_8274, n9251);
  and g17269 (n9252, n_8273, n_8274);
  and g17270 (n9253, n9239, n9252);
  not g17271 (n_8275, n9239);
  not g17272 (n_8276, n9252);
  and g17273 (n9254, n_8275, n_8276);
  not g17274 (n_8277, n9253);
  not g17275 (n_8278, n9254);
  and g17276 (n9255, n_8277, n_8278);
  not g17277 (n_8279, n9192);
  and g17278 (n9256, n_8279, n9255);
  not g17279 (n_8280, n9256);
  and g17280 (n9257, n_8279, n_8280);
  and g17281 (n9258, n9255, n_8280);
  not g17282 (n_8281, n9257);
  not g17283 (n_8282, n9258);
  and g17284 (n9259, n_8281, n_8282);
  not g17285 (n_8283, n9259);
  and g17286 (n9260, n9191, n_8283);
  not g17287 (n_8284, n9191);
  and g17288 (n9261, n_8284, n_8282);
  and g17289 (n9262, n_8281, n9261);
  not g17290 (n_8285, n9260);
  not g17291 (n_8286, n9262);
  and g17292 (n9263, n_8285, n_8286);
  not g17293 (n_8287, n8979);
  and g17294 (n9264, n_8287, n9263);
  not g17295 (n_8288, n9263);
  and g17296 (n9265, n8979, n_8288);
  not g17297 (n_8289, n9264);
  not g17298 (n_8290, n9265);
  and g17299 (n9266, n_8289, n_8290);
  not g17300 (n_8291, n9266);
  and g17301 (n9267, n8978, n_8291);
  not g17302 (n_8292, n8978);
  and g17303 (n9268, n_8292, n_8290);
  and g17304 (n9269, n_8289, n9268);
  not g17305 (n_8293, n9267);
  not g17306 (n_8294, n9269);
  and g17307 (\asquared[63] , n_8293, n_8294);
  not g17308 (n_8295, n9268);
  and g17309 (n9271, n_8289, n_8295);
  and g17310 (n9272, n_8280, n_8285);
  and g17311 (n9273, n_8200, n_8205);
  and g17312 (n9274, n_8248, n_8252);
  and g17313 (n9275, n_8215, n_8219);
  and g17314 (n9276, n9274, n9275);
  not g17315 (n_8296, n9274);
  not g17316 (n_8297, n9275);
  and g17317 (n9277, n_8296, n_8297);
  not g17318 (n_8298, n9276);
  not g17319 (n_8299, n9277);
  and g17320 (n9278, n_8298, n_8299);
  and g17321 (n9279, n_8054, n_8058);
  not g17322 (n_8300, n9278);
  and g17323 (n9280, n_8300, n9279);
  not g17324 (n_8301, n9279);
  and g17325 (n9281, n9278, n_8301);
  not g17326 (n_8302, n9280);
  not g17327 (n_8303, n9281);
  and g17328 (n9282, n_8302, n_8303);
  and g17329 (n9283, n_8036, n_8048);
  and g17330 (n9284, n_8231, n_8235);
  and g17331 (n9285, n9283, n9284);
  not g17332 (n_8304, n9283);
  not g17333 (n_8305, n9284);
  and g17334 (n9286, n_8304, n_8305);
  not g17335 (n_8306, n9285);
  not g17336 (n_8307, n9286);
  and g17337 (n9287, n_8306, n_8307);
  and g17338 (n9288, n_8243, n_8246);
  not g17339 (n_8308, n9287);
  and g17340 (n9289, n_8308, n9288);
  not g17341 (n_8309, n9288);
  and g17342 (n9290, n9287, n_8309);
  not g17343 (n_8310, n9289);
  not g17344 (n_8311, n9290);
  and g17345 (n9291, n_8310, n_8311);
  and g17346 (n9292, n_8191, n_8192);
  not g17347 (n_8312, n9292);
  and g17348 (n9293, n_8197, n_8312);
  not g17349 (n_8313, n9293);
  and g17350 (n9294, n9291, n_8313);
  not g17351 (n_8314, n9291);
  and g17352 (n9295, n_8314, n9293);
  not g17353 (n_8315, n9294);
  not g17354 (n_8316, n9295);
  and g17355 (n9296, n_8315, n_8316);
  and g17356 (n9297, n9072, n9168);
  not g17357 (n_8317, n9072);
  not g17358 (n_8318, n9168);
  and g17359 (n9298, n_8317, n_8318);
  not g17360 (n_8319, n9297);
  not g17361 (n_8320, n9298);
  and g17362 (n9299, n_8319, n_8320);
  not g17363 (n_8321, n9299);
  and g17364 (n9300, n9151, n_8321);
  not g17365 (n_8322, n9151);
  and g17366 (n9301, n_8322, n9299);
  not g17367 (n_8323, n9300);
  not g17368 (n_8324, n9301);
  and g17369 (n9302, n_8323, n_8324);
  and g17370 (n9303, n8993, n9101);
  not g17371 (n_8325, n8993);
  not g17372 (n_8326, n9101);
  and g17373 (n9304, n_8325, n_8326);
  not g17374 (n_8327, n9303);
  not g17375 (n_8328, n9304);
  and g17376 (n9305, n_8327, n_8328);
  not g17377 (n_8329, n9305);
  and g17378 (n9306, n9089, n_8329);
  not g17379 (n_8330, n9089);
  and g17380 (n9307, n_8330, n9305);
  not g17381 (n_8331, n9306);
  not g17382 (n_8332, n9307);
  and g17383 (n9308, n_8331, n_8332);
  and g17384 (n9309, n_8223, n_8227);
  not g17385 (n_8333, n9308);
  and g17386 (n9310, n_8333, n9309);
  not g17387 (n_8334, n9309);
  and g17388 (n9311, n9308, n_8334);
  not g17389 (n_8335, n9310);
  not g17390 (n_8336, n9311);
  and g17391 (n9312, n_8335, n_8336);
  and g17392 (n9313, n9302, n9312);
  not g17393 (n_8337, n9302);
  not g17394 (n_8338, n9312);
  and g17395 (n9314, n_8337, n_8338);
  not g17396 (n_8339, n9313);
  not g17397 (n_8340, n9314);
  and g17398 (n9315, n_8339, n_8340);
  and g17399 (n9316, n9296, n9315);
  not g17400 (n_8341, n9296);
  not g17401 (n_8342, n9315);
  and g17402 (n9317, n_8341, n_8342);
  not g17403 (n_8343, n9316);
  not g17404 (n_8344, n9317);
  and g17405 (n9318, n_8343, n_8344);
  and g17406 (n9319, n9282, n9318);
  not g17407 (n_8345, n9282);
  not g17408 (n_8346, n9318);
  and g17409 (n9320, n_8345, n_8346);
  not g17410 (n_8347, n9273);
  not g17411 (n_8348, n9320);
  and g17412 (n9321, n_8347, n_8348);
  not g17413 (n_8349, n9319);
  and g17414 (n9322, n_8349, n9321);
  not g17415 (n_8350, n9322);
  and g17416 (n9323, n_8347, n_8350);
  and g17417 (n9324, n_8349, n_8350);
  and g17418 (n9325, n_8348, n9324);
  not g17419 (n_8351, n9323);
  not g17420 (n_8352, n9325);
  and g17421 (n9326, n_8351, n_8352);
  and g17422 (n9327, n_8077, n_8211);
  and g17423 (n9328, n9326, n9327);
  not g17424 (n_8353, n9326);
  not g17425 (n_8354, n9327);
  and g17426 (n9329, n_8353, n_8354);
  not g17427 (n_8355, n9328);
  not g17428 (n_8356, n9329);
  and g17429 (n9330, n_8355, n_8356);
  and g17430 (n9331, n_8274, n_8277);
  and g17431 (n9332, n_8266, n_8270);
  and g17432 (n9333, n9055, n9117);
  not g17433 (n_8357, n9055);
  not g17434 (n_8358, n9117);
  and g17435 (n9334, n_8357, n_8358);
  not g17436 (n_8359, n9333);
  not g17437 (n_8360, n9334);
  and g17438 (n9335, n_8359, n_8360);
  not g17439 (n_8361, n9335);
  and g17440 (n9336, n9043, n_8361);
  not g17441 (n_8362, n9043);
  and g17442 (n9337, n_8362, n9335);
  not g17443 (n_8363, n9336);
  not g17444 (n_8364, n9337);
  and g17445 (n9338, n_8363, n_8364);
  and g17446 (n9339, n_8101, n_8116);
  not g17447 (n_8365, n9338);
  and g17448 (n9340, n_8365, n9339);
  not g17449 (n_8366, n9339);
  and g17450 (n9341, n9338, n_8366);
  not g17451 (n_8367, n9340);
  not g17452 (n_8368, n9341);
  and g17453 (n9342, n_8367, n_8368);
  and g17454 (n9343, n_8176, n_8188);
  not g17455 (n_8369, n9342);
  and g17456 (n9344, n_8369, n9343);
  not g17457 (n_8370, n9343);
  and g17458 (n9345, n9342, n_8370);
  not g17459 (n_8371, n9344);
  not g17460 (n_8372, n9345);
  and g17461 (n9346, n_8371, n_8372);
  and g17462 (n9347, n_8062, n_8066);
  and g17463 (n9348, n_8136, n_8151);
  and g17464 (n9349, n9347, n9348);
  not g17465 (n_8373, n9347);
  not g17466 (n_8374, n9348);
  and g17467 (n9350, n_8373, n_8374);
  not g17468 (n_8375, n9349);
  not g17469 (n_8376, n9350);
  and g17470 (n9351, n_8375, n_8376);
  and g17471 (n9352, \a[0] , \a[63] );
  and g17472 (n9353, n9215, n9352);
  not g17473 (n_8378, n9353);
  and g17474 (n9354, n9215, n_8378);
  and g17475 (n9355, n_8238, n9352);
  not g17476 (n_8379, n9354);
  not g17477 (n_8380, n9355);
  and g17478 (n9356, n_8379, n_8380);
  and g17479 (n9357, \a[62] , n2687);
  not g17480 (n_8381, n9357);
  and g17481 (n9358, \a[32] , n_8381);
  and g17482 (n9359, \a[1] , n_8381);
  and g17483 (n9360, \a[62] , n9359);
  not g17484 (n_8382, n9358);
  not g17485 (n_8383, n9360);
  and g17486 (n9361, n_8382, n_8383);
  not g17487 (n_8384, n9356);
  not g17488 (n_8385, n9361);
  and g17489 (n9362, n_8384, n_8385);
  not g17490 (n_8386, n9362);
  and g17491 (n9363, n_8384, n_8386);
  and g17492 (n9364, n_8385, n_8386);
  not g17493 (n_8387, n9363);
  not g17494 (n_8388, n9364);
  and g17495 (n9365, n_8387, n_8388);
  and g17496 (n9366, n2463, n4565);
  and g17497 (n9367, n2301, n5430);
  and g17498 (n9368, n1904, n5083);
  not g17499 (n_8389, n9367);
  not g17500 (n_8390, n9368);
  and g17501 (n9369, n_8389, n_8390);
  not g17502 (n_8391, n9366);
  not g17503 (n_8392, n9369);
  and g17504 (n9370, n_8391, n_8392);
  not g17505 (n_8393, n9370);
  and g17506 (n9371, n_8391, n_8393);
  and g17507 (n9372, \a[25] , \a[38] );
  and g17508 (n9373, \a[26] , \a[37] );
  not g17509 (n_8394, n9372);
  not g17510 (n_8395, n9373);
  and g17511 (n9374, n_8394, n_8395);
  not g17512 (n_8396, n9374);
  and g17513 (n9375, n9371, n_8396);
  and g17514 (n9376, \a[39] , n_8393);
  and g17515 (n9377, \a[24] , n9376);
  not g17516 (n_8397, n9375);
  not g17517 (n_8398, n9377);
  and g17518 (n9378, n_8397, n_8398);
  and g17519 (n9379, n2334, n3319);
  and g17520 (n9380, n2041, n4595);
  and g17521 (n9381, n2331, n3828);
  not g17522 (n_8399, n9380);
  not g17523 (n_8400, n9381);
  and g17524 (n9382, n_8399, n_8400);
  not g17525 (n_8401, n9379);
  not g17526 (n_8402, n9382);
  and g17527 (n9383, n_8401, n_8402);
  not g17528 (n_8403, n9383);
  and g17529 (n9384, \a[36] , n_8403);
  and g17530 (n9385, \a[27] , n9384);
  and g17531 (n9386, \a[28] , \a[35] );
  and g17532 (n9387, \a[29] , \a[34] );
  not g17533 (n_8404, n9386);
  not g17534 (n_8405, n9387);
  and g17535 (n9388, n_8404, n_8405);
  and g17536 (n9389, n_8401, n_8403);
  not g17537 (n_8406, n9388);
  and g17538 (n9390, n_8406, n9389);
  not g17539 (n_8407, n9385);
  not g17540 (n_8408, n9390);
  and g17541 (n9391, n_8407, n_8408);
  not g17542 (n_8409, n9378);
  not g17543 (n_8410, n9391);
  and g17544 (n9392, n_8409, n_8410);
  not g17545 (n_8411, n9392);
  and g17546 (n9393, n_8409, n_8411);
  and g17547 (n9394, n_8410, n_8411);
  not g17548 (n_8412, n9393);
  not g17549 (n_8413, n9394);
  and g17550 (n9395, n_8412, n_8413);
  not g17551 (n_8414, n9365);
  and g17552 (n9396, n_8414, n9395);
  not g17553 (n_8415, n9395);
  and g17554 (n9397, n9365, n_8415);
  not g17555 (n_8416, n9396);
  not g17556 (n_8417, n9397);
  and g17557 (n9398, n_8416, n_8417);
  not g17558 (n_8418, n9398);
  and g17559 (n9399, n9351, n_8418);
  not g17560 (n_8419, n9399);
  and g17561 (n9400, n9351, n_8419);
  and g17562 (n9401, n_8418, n_8419);
  not g17563 (n_8420, n9400);
  not g17564 (n_8421, n9401);
  and g17565 (n9402, n_8420, n_8421);
  not g17566 (n_8422, n9346);
  and g17567 (n9403, n_8422, n9402);
  not g17568 (n_8423, n9402);
  and g17569 (n9404, n9346, n_8423);
  not g17570 (n_8424, n9403);
  not g17571 (n_8425, n9404);
  and g17572 (n9405, n_8424, n_8425);
  not g17573 (n_8426, n9332);
  and g17574 (n9406, n_8426, n9405);
  not g17575 (n_8427, n9405);
  and g17576 (n9407, n9332, n_8427);
  not g17577 (n_8428, n9406);
  not g17578 (n_8429, n9407);
  and g17579 (n9408, n_8428, n_8429);
  not g17580 (n_8430, n9331);
  and g17581 (n9409, n_8430, n9408);
  not g17582 (n_8431, n9408);
  and g17583 (n9410, n9331, n_8431);
  not g17584 (n_8432, n9409);
  not g17585 (n_8433, n9410);
  and g17586 (n9411, n_8432, n_8433);
  and g17587 (n9412, n_8256, n_8262);
  and g17588 (n9413, n_8068, n_8073);
  and g17589 (n9414, \a[46] , \a[54] );
  and g17590 (n9415, n1676, n9414);
  and g17591 (n9416, n6997, n9036);
  and g17592 (n9417, n1052, n5560);
  not g17593 (n_8434, n9416);
  not g17594 (n_8435, n9417);
  and g17595 (n9418, n_8434, n_8435);
  not g17596 (n_8436, n9415);
  not g17597 (n_8437, n9418);
  and g17598 (n9419, n_8436, n_8437);
  not g17599 (n_8438, n9419);
  and g17600 (n9420, n_8436, n_8438);
  and g17601 (n9421, \a[9] , \a[54] );
  and g17602 (n9422, \a[17] , \a[46] );
  not g17603 (n_8439, n9421);
  not g17604 (n_8440, n9422);
  and g17605 (n9423, n_8439, n_8440);
  not g17606 (n_8441, n9423);
  and g17607 (n9424, n9420, n_8441);
  and g17608 (n9425, \a[45] , n_8438);
  and g17609 (n9426, \a[18] , n9425);
  not g17610 (n_8442, n9424);
  not g17611 (n_8443, n9426);
  and g17612 (n9427, n_8442, n_8443);
  and g17613 (n9428, \a[47] , \a[52] );
  and g17614 (n9429, n1843, n9428);
  and g17615 (n9430, n723, n7433);
  and g17616 (n9431, \a[16] , \a[53] );
  and g17617 (n9432, n7730, n9431);
  not g17618 (n_8444, n9430);
  not g17619 (n_8445, n9432);
  and g17620 (n9433, n_8444, n_8445);
  not g17621 (n_8446, n9429);
  not g17622 (n_8447, n9433);
  and g17623 (n9434, n_8446, n_8447);
  not g17624 (n_8448, n9434);
  and g17625 (n9435, \a[53] , n_8448);
  and g17626 (n9436, \a[10] , n9435);
  and g17627 (n9437, \a[11] , \a[52] );
  and g17628 (n9438, \a[16] , \a[47] );
  not g17629 (n_8449, n9437);
  not g17630 (n_8450, n9438);
  and g17631 (n9439, n_8449, n_8450);
  and g17632 (n9440, n_8446, n_8448);
  not g17633 (n_8451, n9439);
  and g17634 (n9441, n_8451, n9440);
  not g17635 (n_8452, n9436);
  not g17636 (n_8453, n9441);
  and g17637 (n9442, n_8452, n_8453);
  not g17638 (n_8454, n9427);
  not g17639 (n_8455, n9442);
  and g17640 (n9443, n_8454, n_8455);
  not g17641 (n_8456, n9443);
  and g17642 (n9444, n_8454, n_8456);
  and g17643 (n9445, n_8455, n_8456);
  not g17644 (n_8457, n9444);
  not g17645 (n_8458, n9445);
  and g17646 (n9446, n_8457, n_8458);
  and g17647 (n9447, n748, n6564);
  and g17648 (n9448, n821, n5888);
  and g17649 (n9449, \a[12] , \a[51] );
  and g17650 (n9450, n7351, n9449);
  not g17651 (n_8459, n9448);
  not g17652 (n_8460, n9450);
  and g17653 (n9451, n_8459, n_8460);
  not g17654 (n_8461, n9447);
  not g17655 (n_8462, n9451);
  and g17656 (n9452, n_8461, n_8462);
  not g17657 (n_8463, n9452);
  and g17658 (n9453, n7351, n_8463);
  and g17659 (n9454, n_8461, n_8463);
  and g17660 (n9455, \a[13] , \a[50] );
  not g17661 (n_8464, n9449);
  not g17662 (n_8465, n9455);
  and g17663 (n9456, n_8464, n_8465);
  not g17664 (n_8466, n9456);
  and g17665 (n9457, n9454, n_8466);
  not g17666 (n_8467, n9453);
  not g17667 (n_8468, n9457);
  and g17668 (n9458, n_8467, n_8468);
  not g17669 (n_8469, n9446);
  not g17670 (n_8470, n9458);
  and g17671 (n9459, n_8469, n_8470);
  not g17672 (n_8471, n9459);
  and g17673 (n9460, n_8469, n_8471);
  and g17674 (n9461, n_8470, n_8471);
  not g17675 (n_8472, n9460);
  not g17676 (n_8473, n9461);
  and g17677 (n9462, n_8472, n_8473);
  and g17678 (n9463, \a[6] , \a[57] );
  and g17679 (n9464, \a[20] , \a[43] );
  not g17680 (n_8474, n9463);
  not g17681 (n_8475, n9464);
  and g17682 (n9465, n_8474, n_8475);
  and g17683 (n9466, n9463, n9464);
  not g17684 (n_8476, n9466);
  not g17687 (n_8477, n9465);
  not g17689 (n_8478, n9469);
  and g17690 (n9470, n_8476, n_8478);
  and g17691 (n9471, n_8477, n9470);
  and g17692 (n9472, \a[40] , n_8478);
  and g17693 (n9473, \a[23] , n9472);
  not g17694 (n_8479, n9471);
  not g17695 (n_8480, n9473);
  and g17696 (n9474, n_8479, n_8480);
  and g17697 (n9475, \a[30] , \a[33] );
  not g17698 (n_8481, n3812);
  not g17699 (n_8482, n9475);
  and g17700 (n9476, n_8481, n_8482);
  and g17701 (n9477, n3812, n9475);
  not g17702 (n_8483, n9477);
  not g17705 (n_8484, n9476);
  not g17707 (n_8485, n9480);
  and g17708 (n9481, \a[49] , n_8485);
  and g17709 (n9482, \a[14] , n9481);
  and g17710 (n9483, n_8483, n_8485);
  and g17711 (n9484, n_8484, n9483);
  not g17712 (n_8486, n9482);
  not g17713 (n_8487, n9484);
  and g17714 (n9485, n_8486, n_8487);
  not g17715 (n_8488, n9474);
  not g17716 (n_8489, n9485);
  and g17717 (n9486, n_8488, n_8489);
  not g17718 (n_8490, n9486);
  and g17719 (n9487, n_8488, n_8490);
  and g17720 (n9488, n_8489, n_8490);
  not g17721 (n_8491, n9487);
  not g17722 (n_8492, n9488);
  and g17723 (n9489, n_8491, n_8492);
  and g17724 (n9490, \a[44] , \a[55] );
  and g17725 (n9491, n1856, n9490);
  and g17726 (n9492, n380, n9161);
  and g17727 (n9493, \a[44] , \a[56] );
  and g17728 (n9494, n1662, n9493);
  not g17729 (n_8493, n9492);
  not g17730 (n_8494, n9494);
  and g17731 (n9495, n_8493, n_8494);
  not g17732 (n_8495, n9491);
  not g17733 (n_8496, n9495);
  and g17734 (n9496, n_8495, n_8496);
  not g17735 (n_8497, n9496);
  and g17736 (n9497, \a[56] , n_8497);
  and g17737 (n9498, \a[7] , n9497);
  and g17738 (n9499, \a[8] , \a[55] );
  and g17739 (n9500, \a[19] , \a[44] );
  not g17740 (n_8498, n9499);
  not g17741 (n_8499, n9500);
  and g17742 (n9501, n_8498, n_8499);
  and g17743 (n9502, n_8495, n_8497);
  not g17744 (n_8500, n9501);
  and g17745 (n9503, n_8500, n9502);
  not g17746 (n_8501, n9498);
  not g17747 (n_8502, n9503);
  and g17748 (n9504, n_8501, n_8502);
  not g17749 (n_8503, n9489);
  not g17750 (n_8504, n9504);
  and g17751 (n9505, n_8503, n_8504);
  not g17752 (n_8505, n9505);
  and g17753 (n9506, n_8503, n_8505);
  and g17754 (n9507, n_8504, n_8505);
  not g17755 (n_8506, n9506);
  not g17756 (n_8507, n9507);
  and g17757 (n9508, n_8506, n_8507);
  and g17758 (n9509, \a[59] , \a[60] );
  and g17759 (n9510, n209, n9509);
  and g17760 (n9511, n252, n8905);
  and g17761 (n9512, \a[60] , \a[61] );
  and g17762 (n9513, n218, n9512);
  not g17763 (n_8508, n9511);
  not g17764 (n_8509, n9513);
  and g17765 (n9514, n_8508, n_8509);
  not g17766 (n_8510, n9510);
  not g17767 (n_8511, n9514);
  and g17768 (n9515, n_8510, n_8511);
  not g17769 (n_8512, n9515);
  and g17770 (n9516, \a[2] , n_8512);
  and g17771 (n9517, \a[61] , n9516);
  and g17772 (n9518, n_8510, n_8512);
  and g17773 (n9519, \a[3] , \a[60] );
  and g17774 (n9520, \a[4] , \a[59] );
  not g17775 (n_8513, n9519);
  not g17776 (n_8514, n9520);
  and g17777 (n9521, n_8513, n_8514);
  not g17778 (n_8515, n9521);
  and g17779 (n9522, n9518, n_8515);
  not g17780 (n_8516, n9517);
  not g17781 (n_8517, n9522);
  and g17782 (n9523, n_8516, n_8517);
  not g17783 (n_8518, n9523);
  and g17784 (n9524, n9133, n_8518);
  not g17785 (n_8519, n9133);
  and g17786 (n9525, n_8519, n9523);
  not g17787 (n_8520, n9524);
  not g17788 (n_8521, n9525);
  and g17789 (n9526, n_8520, n_8521);
  and g17790 (n9527, \a[21] , \a[42] );
  and g17791 (n9528, \a[22] , \a[41] );
  not g17792 (n_8522, n9527);
  not g17793 (n_8523, n9528);
  and g17794 (n9529, n_8522, n_8523);
  and g17795 (n9530, n1574, n5344);
  not g17796 (n_8524, n9530);
  not g17799 (n_8525, n9529);
  not g17801 (n_8526, n9533);
  and g17802 (n9534, \a[58] , n_8526);
  and g17803 (n9535, \a[5] , n9534);
  and g17804 (n9536, n_8524, n_8526);
  and g17805 (n9537, n_8525, n9536);
  not g17806 (n_8527, n9535);
  not g17807 (n_8528, n9537);
  and g17808 (n9538, n_8527, n_8528);
  not g17809 (n_8529, n9526);
  not g17810 (n_8530, n9538);
  and g17811 (n9539, n_8529, n_8530);
  and g17812 (n9540, n9526, n9538);
  not g17813 (n_8531, n9539);
  not g17814 (n_8532, n9540);
  and g17815 (n9541, n_8531, n_8532);
  and g17816 (n9542, n9508, n9541);
  not g17817 (n_8533, n9508);
  not g17818 (n_8534, n9541);
  and g17819 (n9543, n_8533, n_8534);
  not g17820 (n_8535, n9542);
  not g17821 (n_8536, n9543);
  and g17822 (n9544, n_8535, n_8536);
  not g17823 (n_8537, n9462);
  not g17824 (n_8538, n9544);
  and g17825 (n9545, n_8537, n_8538);
  and g17826 (n9546, n9462, n9544);
  not g17827 (n_8539, n9545);
  not g17828 (n_8540, n9546);
  and g17829 (n9547, n_8539, n_8540);
  not g17830 (n_8541, n9413);
  and g17831 (n9548, n_8541, n9547);
  not g17832 (n_8542, n9548);
  and g17833 (n9549, n_8541, n_8542);
  and g17834 (n9550, n9547, n_8542);
  not g17835 (n_8543, n9549);
  not g17836 (n_8544, n9550);
  and g17837 (n9551, n_8543, n_8544);
  not g17838 (n_8545, n9412);
  not g17839 (n_8546, n9551);
  and g17840 (n9552, n_8545, n_8546);
  not g17841 (n_8547, n9552);
  and g17842 (n9553, n_8545, n_8547);
  and g17843 (n9554, n_8546, n_8547);
  not g17844 (n_8548, n9553);
  not g17845 (n_8549, n9554);
  and g17846 (n9555, n_8548, n_8549);
  not g17847 (n_8550, n9555);
  and g17848 (n9556, n9411, n_8550);
  not g17849 (n_8551, n9556);
  and g17850 (n9557, n9411, n_8551);
  and g17851 (n9558, n_8550, n_8551);
  not g17852 (n_8552, n9557);
  not g17853 (n_8553, n9558);
  and g17854 (n9559, n_8552, n_8553);
  not g17855 (n_8554, n9330);
  and g17856 (n9560, n_8554, n9559);
  not g17857 (n_8555, n9559);
  and g17858 (n9561, n9330, n_8555);
  not g17859 (n_8556, n9560);
  not g17860 (n_8557, n9561);
  and g17861 (n9562, n_8556, n_8557);
  not g17862 (n_8558, n9562);
  and g17863 (n9563, n9272, n_8558);
  not g17864 (n_8559, n9272);
  and g17865 (n9564, n_8559, n9562);
  not g17866 (n_8560, n9563);
  not g17867 (n_8561, n9564);
  and g17868 (n9565, n_8560, n_8561);
  not g17869 (n_8562, n9271);
  not g17870 (n_8563, n9565);
  and g17871 (n9566, n_8562, n_8563);
  and g17872 (n9567, n9271, n9565);
  or g17873 (\asquared[64] , n9566, n9567);
  and g17874 (n9569, n_8562, n_8560);
  not g17875 (n_8564, n9569);
  and g17876 (n9570, n_8561, n_8564);
  and g17877 (n9571, n_8432, n_8551);
  and g17878 (n9572, n_8542, n_8547);
  and g17879 (n9573, n_8425, n_8428);
  and g17880 (n9574, n_8533, n9541);
  not g17881 (n_8565, n9574);
  and g17882 (n9575, n_8539, n_8565);
  and g17883 (n9576, n_8376, n_8419);
  and g17884 (n9577, n9575, n9576);
  not g17885 (n_8566, n9575);
  not g17886 (n_8567, n9576);
  and g17887 (n9578, n_8566, n_8567);
  not g17888 (n_8568, n9577);
  not g17889 (n_8569, n9578);
  and g17890 (n9579, n_8568, n_8569);
  and g17891 (n9580, n_8414, n_8415);
  not g17892 (n_8570, n9580);
  and g17893 (n9581, n_8411, n_8570);
  and g17894 (n9582, n9420, n9470);
  not g17895 (n_8571, n9420);
  not g17896 (n_8572, n9470);
  and g17897 (n9583, n_8571, n_8572);
  not g17898 (n_8573, n9582);
  not g17899 (n_8574, n9583);
  and g17900 (n9584, n_8573, n_8574);
  not g17901 (n_8575, n9584);
  and g17902 (n9585, n9389, n_8575);
  not g17903 (n_8576, n9389);
  and g17904 (n9586, n_8576, n9584);
  not g17905 (n_8577, n9585);
  not g17906 (n_8578, n9586);
  and g17907 (n9587, n_8577, n_8578);
  and g17908 (n9588, n9518, n9536);
  not g17909 (n_8579, n9518);
  not g17910 (n_8580, n9536);
  and g17911 (n9589, n_8579, n_8580);
  not g17912 (n_8581, n9588);
  not g17913 (n_8582, n9589);
  and g17914 (n9590, n_8581, n_8582);
  not g17915 (n_8583, n9590);
  and g17916 (n9591, n9502, n_8583);
  not g17917 (n_8584, n9502);
  and g17918 (n9592, n_8584, n9590);
  not g17919 (n_8585, n9591);
  not g17920 (n_8586, n9592);
  and g17921 (n9593, n_8585, n_8586);
  not g17922 (n_8587, n9587);
  not g17923 (n_8588, n9593);
  and g17924 (n9594, n_8587, n_8588);
  and g17925 (n9595, n9587, n9593);
  not g17926 (n_8589, n9594);
  not g17927 (n_8590, n9595);
  and g17928 (n9596, n_8589, n_8590);
  not g17929 (n_8591, n9581);
  and g17930 (n9597, n_8591, n9596);
  not g17931 (n_8592, n9596);
  and g17932 (n9598, n9581, n_8592);
  not g17933 (n_8593, n9597);
  not g17934 (n_8594, n9598);
  and g17935 (n9599, n_8593, n_8594);
  not g17936 (n_8595, n9579);
  not g17937 (n_8596, n9599);
  and g17938 (n9600, n_8595, n_8596);
  and g17939 (n9601, n9579, n9599);
  not g17940 (n_8597, n9600);
  not g17941 (n_8598, n9601);
  and g17942 (n9602, n_8597, n_8598);
  not g17943 (n_8599, n9573);
  and g17944 (n9603, n_8599, n9602);
  not g17945 (n_8600, n9603);
  and g17946 (n9604, n_8599, n_8600);
  and g17947 (n9605, n9602, n_8600);
  not g17948 (n_8601, n9604);
  not g17949 (n_8602, n9605);
  and g17950 (n9606, n_8601, n_8602);
  not g17951 (n_8603, n9572);
  not g17952 (n_8604, n9606);
  and g17953 (n9607, n_8603, n_8604);
  not g17954 (n_8605, n9607);
  and g17955 (n9608, n_8603, n_8605);
  and g17956 (n9609, n_8604, n_8605);
  not g17957 (n_8606, n9608);
  not g17958 (n_8607, n9609);
  and g17959 (n9610, n_8606, n_8607);
  not g17960 (n_8608, n9571);
  not g17961 (n_8609, n9610);
  and g17962 (n9611, n_8608, n_8609);
  not g17963 (n_8610, n9611);
  and g17964 (n9612, n_8608, n_8610);
  and g17965 (n9613, n_8609, n_8610);
  not g17966 (n_8611, n9612);
  not g17967 (n_8612, n9613);
  and g17968 (n9614, n_8611, n_8612);
  and g17969 (n9615, n_8315, n_8343);
  and g17970 (n9616, \a[7] , \a[57] );
  not g17971 (n_8613, n5899);
  not g17972 (n_8614, n9616);
  and g17973 (n9617, n_8613, n_8614);
  and g17974 (n9618, \a[17] , \a[57] );
  and g17975 (n9619, n6980, n9618);
  and g17976 (n9620, \a[58] , n6610);
  and g17977 (n9621, \a[17] , n9620);
  and g17978 (n9622, n335, n8436);
  not g17979 (n_8615, n9621);
  not g17980 (n_8616, n9622);
  and g17981 (n9623, n_8615, n_8616);
  not g17982 (n_8617, n9619);
  not g17983 (n_8618, n9623);
  and g17984 (n9624, n_8617, n_8618);
  not g17985 (n_8619, n9624);
  and g17986 (n9625, n_8617, n_8619);
  not g17987 (n_8620, n9617);
  and g17988 (n9626, n_8620, n9625);
  and g17989 (n9627, \a[58] , n_8619);
  and g17990 (n9628, \a[6] , n9627);
  not g17991 (n_8621, n9626);
  not g17992 (n_8622, n9628);
  and g17993 (n9629, n_8621, n_8622);
  and g17994 (n9630, n1574, n5018);
  and g17995 (n9631, n1693, n4639);
  and g17996 (n9632, n1494, n5296);
  not g17997 (n_8623, n9631);
  not g17998 (n_8624, n9632);
  and g17999 (n9633, n_8623, n_8624);
  not g18000 (n_8625, n9630);
  not g18001 (n_8626, n9633);
  and g18002 (n9634, n_8625, n_8626);
  not g18003 (n_8627, n9634);
  and g18004 (n9635, \a[44] , n_8627);
  and g18005 (n9636, \a[20] , n9635);
  and g18006 (n9637, n_8625, n_8627);
  and g18007 (n9638, \a[21] , \a[43] );
  and g18008 (n9639, \a[22] , \a[42] );
  not g18009 (n_8628, n9638);
  not g18010 (n_8629, n9639);
  and g18011 (n9640, n_8628, n_8629);
  not g18012 (n_8630, n9640);
  and g18013 (n9641, n9637, n_8630);
  not g18014 (n_8631, n9636);
  not g18015 (n_8632, n9641);
  and g18016 (n9642, n_8631, n_8632);
  not g18017 (n_8633, n9629);
  not g18018 (n_8634, n9642);
  and g18019 (n9643, n_8633, n_8634);
  not g18020 (n_8635, n9643);
  and g18021 (n9644, n_8633, n_8635);
  and g18022 (n9645, n_8634, n_8635);
  not g18023 (n_8636, n9644);
  not g18024 (n_8637, n9645);
  and g18025 (n9646, n_8636, n_8637);
  and g18026 (n9647, n1904, n4171);
  and g18027 (n9648, n1547, n3984);
  and g18028 (n9649, n1666, n5413);
  not g18029 (n_8638, n9648);
  not g18030 (n_8639, n9649);
  and g18031 (n9650, n_8638, n_8639);
  not g18032 (n_8640, n9647);
  not g18033 (n_8641, n9650);
  and g18034 (n9651, n_8640, n_8641);
  not g18035 (n_8642, n9651);
  and g18036 (n9652, \a[41] , n_8642);
  and g18037 (n9653, \a[23] , n9652);
  and g18038 (n9654, n_8640, n_8642);
  and g18039 (n9655, \a[24] , \a[40] );
  and g18040 (n9656, \a[25] , \a[39] );
  not g18041 (n_8643, n9655);
  not g18042 (n_8644, n9656);
  and g18043 (n9657, n_8643, n_8644);
  not g18044 (n_8645, n9657);
  and g18045 (n9658, n9654, n_8645);
  not g18046 (n_8646, n9653);
  not g18047 (n_8647, n9658);
  and g18048 (n9659, n_8646, n_8647);
  not g18049 (n_8648, n9646);
  not g18050 (n_8649, n9659);
  and g18051 (n9660, n_8648, n_8649);
  not g18052 (n_8650, n9660);
  and g18053 (n9661, n_8648, n_8650);
  and g18054 (n9662, n_8649, n_8650);
  not g18055 (n_8651, n9661);
  not g18056 (n_8652, n9662);
  and g18057 (n9663, n_8651, n_8652);
  and g18058 (n9664, \a[8] , \a[56] );
  not g18059 (n_8653, n6642);
  not g18060 (n_8654, n9664);
  and g18061 (n9665, n_8653, n_8654);
  and g18062 (n9666, \a[48] , \a[56] );
  and g18063 (n9667, n1509, n9666);
  not g18064 (n_8655, n9667);
  not g18067 (n_8656, n9665);
  not g18069 (n_8657, n9670);
  and g18070 (n9671, n_8655, n_8657);
  and g18071 (n9672, n_8656, n9671);
  and g18072 (n9673, \a[38] , n_8657);
  and g18073 (n9674, \a[26] , n9673);
  not g18074 (n_8658, n9672);
  not g18075 (n_8659, n9674);
  and g18076 (n9675, n_8658, n_8659);
  and g18077 (n9676, n2334, n3828);
  and g18078 (n9677, n2041, n5031);
  and g18079 (n9678, n2331, n3687);
  not g18080 (n_8660, n9677);
  not g18081 (n_8661, n9678);
  and g18082 (n9679, n_8660, n_8661);
  not g18083 (n_8662, n9676);
  not g18084 (n_8663, n9679);
  and g18085 (n9680, n_8662, n_8663);
  not g18086 (n_8664, n9680);
  and g18087 (n9681, n4059, n_8664);
  and g18088 (n9682, n_8662, n_8664);
  and g18089 (n9683, \a[28] , \a[36] );
  and g18090 (n9684, \a[29] , \a[35] );
  not g18091 (n_8665, n9683);
  not g18092 (n_8666, n9684);
  and g18093 (n9685, n_8665, n_8666);
  not g18094 (n_8667, n9685);
  and g18095 (n9686, n9682, n_8667);
  not g18096 (n_8668, n9681);
  not g18097 (n_8669, n9686);
  and g18098 (n9687, n_8668, n_8669);
  not g18099 (n_8670, n9675);
  not g18100 (n_8671, n9687);
  and g18101 (n9688, n_8670, n_8671);
  not g18102 (n_8672, n9688);
  and g18103 (n9689, n_8670, n_8672);
  and g18104 (n9690, n_8671, n_8672);
  not g18105 (n_8673, n9689);
  not g18106 (n_8674, n9690);
  and g18107 (n9691, n_8673, n_8674);
  and g18108 (n9692, \a[30] , \a[34] );
  not g18109 (n_8675, n2598);
  not g18110 (n_8676, n9692);
  and g18111 (n9693, n_8675, n_8676);
  and g18112 (n9694, n2865, n4150);
  not g18113 (n_8677, n9694);
  and g18114 (n9695, n8868, n_8677);
  not g18115 (n_8678, n9693);
  and g18116 (n9696, n_8678, n9695);
  not g18117 (n_8679, n9696);
  and g18118 (n9697, n8868, n_8679);
  and g18119 (n9698, n_8677, n_8679);
  and g18120 (n9699, n_8678, n9698);
  not g18121 (n_8680, n9697);
  not g18122 (n_8681, n9699);
  and g18123 (n9700, n_8680, n_8681);
  not g18124 (n_8682, n9691);
  not g18125 (n_8683, n9700);
  and g18126 (n9701, n_8682, n_8683);
  not g18127 (n_8684, n9701);
  and g18128 (n9702, n_8682, n_8684);
  and g18129 (n9703, n_8683, n_8684);
  not g18130 (n_8685, n9702);
  not g18131 (n_8686, n9703);
  and g18132 (n9704, n_8685, n_8686);
  and g18133 (n9705, n1149, n5560);
  and g18134 (n9706, \a[18] , \a[46] );
  and g18135 (n9707, \a[19] , \a[45] );
  not g18136 (n_8687, n9706);
  not g18137 (n_8688, n9707);
  and g18138 (n9708, n_8687, n_8688);
  not g18139 (n_8689, n9705);
  not g18140 (n_8690, n9708);
  and g18141 (n9709, n_8689, n_8690);
  and g18142 (n9710, n8903, n9709);
  not g18143 (n_8691, n9710);
  and g18144 (n9711, n8903, n_8691);
  and g18145 (n9712, n_8689, n_8691);
  and g18146 (n9713, n_8690, n9712);
  not g18147 (n_8692, n9711);
  not g18148 (n_8693, n9713);
  and g18149 (n9714, n_8692, n_8693);
  and g18150 (n9715, n_8378, n_8386);
  not g18151 (n_8694, n9714);
  and g18152 (n9716, n_8694, n9715);
  not g18153 (n_8695, n9715);
  and g18154 (n9717, n9714, n_8695);
  not g18155 (n_8696, n9716);
  not g18156 (n_8697, n9717);
  and g18157 (n9718, n_8696, n_8697);
  and g18158 (n9719, n209, n9512);
  and g18159 (n9720, n252, n9085);
  and g18160 (n9721, \a[61] , \a[62] );
  and g18161 (n9722, n218, n9721);
  not g18162 (n_8698, n9720);
  not g18163 (n_8699, n9722);
  and g18164 (n9723, n_8698, n_8699);
  not g18165 (n_8700, n9719);
  not g18166 (n_8701, n9723);
  and g18167 (n9724, n_8700, n_8701);
  not g18168 (n_8702, n9724);
  and g18169 (n9725, \a[62] , n_8702);
  and g18170 (n9726, \a[2] , n9725);
  and g18171 (n9727, n_8700, n_8702);
  and g18172 (n9728, \a[3] , \a[61] );
  and g18173 (n9729, \a[4] , \a[60] );
  not g18174 (n_8703, n9728);
  not g18175 (n_8704, n9729);
  and g18176 (n9730, n_8703, n_8704);
  not g18177 (n_8705, n9730);
  and g18178 (n9731, n9727, n_8705);
  not g18179 (n_8706, n9726);
  not g18180 (n_8707, n9731);
  and g18181 (n9732, n_8706, n_8707);
  not g18182 (n_8708, n9718);
  not g18183 (n_8709, n9732);
  and g18184 (n9733, n_8708, n_8709);
  and g18185 (n9734, n9718, n9732);
  not g18186 (n_8710, n9733);
  not g18187 (n_8711, n9734);
  and g18188 (n9735, n_8710, n_8711);
  and g18189 (n9736, n9704, n9735);
  not g18190 (n_8712, n9704);
  not g18191 (n_8713, n9735);
  and g18192 (n9737, n_8712, n_8713);
  not g18193 (n_8714, n9736);
  not g18194 (n_8715, n9737);
  and g18195 (n9738, n_8714, n_8715);
  not g18196 (n_8716, n9663);
  not g18197 (n_8717, n9738);
  and g18198 (n9739, n_8716, n_8717);
  and g18199 (n9740, n9663, n9738);
  not g18200 (n_8718, n9739);
  not g18201 (n_8719, n9740);
  and g18202 (n9741, n_8718, n_8719);
  not g18203 (n_8720, n9615);
  and g18204 (n9742, n_8720, n9741);
  not g18205 (n_8721, n9741);
  and g18206 (n9743, n9615, n_8721);
  not g18207 (n_8722, n9742);
  not g18208 (n_8723, n9743);
  and g18209 (n9744, n_8722, n_8723);
  and g18210 (n9745, n_8320, n_8324);
  and g18211 (n9746, n_8360, n_8364);
  and g18212 (n9747, n9745, n9746);
  not g18213 (n_8724, n9745);
  not g18214 (n_8725, n9746);
  and g18215 (n9748, n_8724, n_8725);
  not g18216 (n_8726, n9747);
  not g18217 (n_8727, n9748);
  and g18218 (n9749, n_8726, n_8727);
  and g18219 (n9750, n_8328, n_8332);
  not g18220 (n_8728, n9749);
  and g18221 (n9751, n_8728, n9750);
  not g18222 (n_8729, n9750);
  and g18223 (n9752, n9749, n_8729);
  not g18224 (n_8730, n9751);
  not g18225 (n_8731, n9752);
  and g18226 (n9753, n_8730, n_8731);
  and g18227 (n9754, n_8368, n_8372);
  and g18228 (n9755, n_8336, n_8339);
  not g18229 (n_8732, n9754);
  not g18230 (n_8733, n9755);
  and g18231 (n9756, n_8732, n_8733);
  not g18232 (n_8734, n9756);
  and g18233 (n9757, n_8732, n_8734);
  and g18234 (n9758, n_8733, n_8734);
  not g18235 (n_8735, n9757);
  not g18236 (n_8736, n9758);
  and g18237 (n9759, n_8735, n_8736);
  not g18238 (n_8737, n9759);
  and g18239 (n9760, n9753, n_8737);
  not g18240 (n_8738, n9753);
  and g18241 (n9761, n_8738, n9759);
  not g18242 (n_8739, n9761);
  and g18243 (n9762, n9744, n_8739);
  not g18244 (n_8740, n9760);
  and g18245 (n9763, n_8740, n9762);
  not g18246 (n_8741, n9763);
  and g18247 (n9764, n9744, n_8741);
  and g18248 (n9765, n_8739, n_8741);
  and g18249 (n9766, n_8740, n9765);
  not g18250 (n_8742, n9764);
  not g18251 (n_8743, n9766);
  and g18252 (n9767, n_8742, n_8743);
  and g18253 (n9768, n9371, n9454);
  not g18254 (n_8744, n9371);
  not g18255 (n_8745, n9454);
  and g18256 (n9769, n_8744, n_8745);
  not g18257 (n_8746, n9768);
  not g18258 (n_8747, n9769);
  and g18259 (n9770, n_8746, n_8747);
  not g18260 (n_8748, n9770);
  and g18261 (n9771, n9440, n_8748);
  not g18262 (n_8749, n9440);
  and g18263 (n9772, n_8749, n9770);
  not g18264 (n_8750, n9771);
  not g18265 (n_8751, n9772);
  and g18266 (n9773, n_8750, n_8751);
  and g18267 (n9774, n_8490, n_8505);
  not g18268 (n_8752, n9773);
  and g18269 (n9775, n_8752, n9774);
  not g18270 (n_8753, n9774);
  and g18271 (n9776, n9773, n_8753);
  not g18272 (n_8754, n9775);
  not g18273 (n_8755, n9776);
  and g18274 (n9777, n_8754, n_8755);
  and g18275 (n9778, n_8456, n_8471);
  not g18276 (n_8756, n9777);
  and g18277 (n9779, n_8756, n9778);
  not g18278 (n_8757, n9778);
  and g18279 (n9780, n9777, n_8757);
  not g18280 (n_8758, n9779);
  not g18281 (n_8759, n9780);
  and g18282 (n9781, n_8758, n_8759);
  and g18283 (n9782, n_8299, n_8303);
  not g18284 (n_8760, n9781);
  and g18285 (n9783, n_8760, n9782);
  not g18286 (n_8761, n9782);
  and g18287 (n9784, n9781, n_8761);
  not g18288 (n_8762, n9783);
  not g18289 (n_8763, n9784);
  and g18290 (n9785, n_8762, n_8763);
  and g18291 (n9786, n_8307, n_8311);
  and g18292 (n9787, n_8519, n_8518);
  not g18293 (n_8764, n9787);
  and g18294 (n9788, n_8531, n_8764);
  and g18295 (n9789, n9786, n9788);
  not g18296 (n_8765, n9786);
  not g18297 (n_8766, n9788);
  and g18298 (n9790, n_8765, n_8766);
  not g18299 (n_8767, n9789);
  not g18300 (n_8768, n9790);
  and g18301 (n9791, n_8767, n_8768);
  and g18302 (n9792, \a[62] , \a[63] );
  and g18303 (n9793, n2687, n9792);
  not g18304 (n_8769, n9793);
  and g18305 (n9794, n9357, n_8769);
  and g18306 (n9795, \a[63] , n9359);
  not g18307 (n_8770, n9794);
  not g18308 (n_8771, n9795);
  and g18309 (n9796, n_8770, n_8771);
  not g18310 (n_8772, n9483);
  not g18311 (n_8773, n9796);
  and g18312 (n9797, n_8772, n_8773);
  not g18313 (n_8774, n9797);
  and g18314 (n9798, n_8772, n_8774);
  and g18315 (n9799, n_8773, n_8774);
  not g18316 (n_8775, n9798);
  not g18317 (n_8776, n9799);
  and g18318 (n9800, n_8775, n_8776);
  and g18319 (n9801, \a[49] , \a[55] );
  and g18320 (n9802, n1517, n9801);
  and g18321 (n9803, n484, n7701);
  not g18322 (n_8777, n9802);
  not g18323 (n_8778, n9803);
  and g18324 (n9804, n_8777, n_8778);
  and g18325 (n9805, \a[10] , \a[54] );
  and g18326 (n9806, \a[15] , \a[49] );
  and g18327 (n9807, n9805, n9806);
  not g18328 (n_8779, n9804);
  not g18329 (n_8780, n9807);
  and g18330 (n9808, n_8779, n_8780);
  not g18331 (n_8781, n9808);
  and g18332 (n9809, n_8780, n_8781);
  not g18333 (n_8782, n9805);
  not g18334 (n_8783, n9806);
  and g18335 (n9810, n_8782, n_8783);
  not g18336 (n_8784, n9810);
  and g18337 (n9811, n9809, n_8784);
  and g18338 (n9812, \a[55] , n_8781);
  and g18339 (n9813, \a[9] , n9812);
  not g18340 (n_8785, n9811);
  not g18341 (n_8786, n9813);
  and g18342 (n9814, n_8785, n_8786);
  and g18343 (n9815, n602, n7433);
  and g18344 (n9816, n818, n7232);
  and g18345 (n9817, n748, n6968);
  not g18346 (n_8787, n9816);
  not g18347 (n_8788, n9817);
  and g18348 (n9818, n_8787, n_8788);
  not g18349 (n_8789, n9815);
  not g18350 (n_8790, n9818);
  and g18351 (n9819, n_8789, n_8790);
  not g18352 (n_8791, n9819);
  and g18353 (n9820, \a[51] , n_8791);
  and g18354 (n9821, \a[13] , n9820);
  and g18355 (n9822, \a[11] , \a[53] );
  and g18356 (n9823, \a[12] , \a[52] );
  not g18357 (n_8792, n9822);
  not g18358 (n_8793, n9823);
  and g18359 (n9824, n_8792, n_8793);
  and g18360 (n9825, n_8789, n_8791);
  not g18361 (n_8794, n9824);
  and g18362 (n9826, n_8794, n9825);
  not g18363 (n_8795, n9821);
  not g18364 (n_8796, n9826);
  and g18365 (n9827, n_8795, n_8796);
  not g18366 (n_8797, n9814);
  not g18367 (n_8798, n9827);
  and g18368 (n9828, n_8797, n_8798);
  not g18369 (n_8799, n9828);
  and g18370 (n9829, n_8797, n_8799);
  and g18371 (n9830, n_8798, n_8799);
  not g18372 (n_8800, n9829);
  not g18373 (n_8801, n9830);
  and g18374 (n9831, n_8800, n_8801);
  not g18375 (n_8802, n9800);
  and g18376 (n9832, n_8802, n9831);
  not g18377 (n_8803, n9831);
  and g18378 (n9833, n9800, n_8803);
  not g18379 (n_8804, n9832);
  not g18380 (n_8805, n9833);
  and g18381 (n9834, n_8804, n_8805);
  not g18382 (n_8806, n9834);
  and g18383 (n9835, n9791, n_8806);
  not g18384 (n_8807, n9835);
  and g18385 (n9836, n9791, n_8807);
  and g18386 (n9837, n_8806, n_8807);
  not g18387 (n_8808, n9836);
  not g18388 (n_8809, n9837);
  and g18389 (n9838, n_8808, n_8809);
  not g18390 (n_8810, n9785);
  and g18391 (n9839, n_8810, n9838);
  not g18392 (n_8811, n9838);
  and g18393 (n9840, n9785, n_8811);
  not g18394 (n_8812, n9839);
  not g18395 (n_8813, n9840);
  and g18396 (n9841, n_8812, n_8813);
  not g18397 (n_8814, n9324);
  and g18398 (n9842, n_8814, n9841);
  not g18399 (n_8815, n9841);
  and g18400 (n9843, n9324, n_8815);
  not g18401 (n_8816, n9842);
  not g18402 (n_8817, n9843);
  and g18403 (n9844, n_8816, n_8817);
  not g18404 (n_8818, n9767);
  and g18405 (n9845, n_8818, n9844);
  not g18406 (n_8819, n9844);
  and g18407 (n9846, n9767, n_8819);
  not g18408 (n_8820, n9845);
  not g18409 (n_8821, n9846);
  and g18410 (n9847, n_8820, n_8821);
  not g18411 (n_8822, n9614);
  and g18412 (n9848, n_8822, n9847);
  not g18413 (n_8823, n9847);
  and g18414 (n9849, n9614, n_8823);
  not g18415 (n_8824, n9848);
  not g18416 (n_8825, n9849);
  and g18417 (n9850, n_8824, n_8825);
  and g18418 (n9851, n_8356, n_8557);
  not g18419 (n_8826, n9850);
  and g18420 (n9852, n_8826, n9851);
  not g18421 (n_8827, n9851);
  and g18422 (n9853, n9850, n_8827);
  not g18423 (n_8828, n9852);
  not g18424 (n_8829, n9853);
  and g18425 (n9854, n_8828, n_8829);
  not g18426 (n_8830, n9854);
  and g18427 (n9855, n9570, n_8830);
  not g18428 (n_8831, n9570);
  and g18429 (n9856, n_8831, n_8828);
  and g18430 (n9857, n_8829, n9856);
  not g18431 (n_8832, n9855);
  not g18432 (n_8833, n9857);
  and g18433 (\asquared[65] , n_8832, n_8833);
  not g18434 (n_8834, n9856);
  and g18435 (n9859, n_8829, n_8834);
  and g18436 (n9860, n_8610, n_8824);
  and g18437 (n9861, n_8816, n_8820);
  and g18438 (n9862, n_8722, n_8741);
  and g18439 (n9863, n_8763, n_8813);
  and g18440 (n9864, n_8712, n9735);
  not g18441 (n_8835, n9864);
  and g18442 (n9865, n_8718, n_8835);
  and g18443 (n9866, n_8768, n_8807);
  and g18444 (n9867, n9865, n9866);
  not g18445 (n_8836, n9865);
  not g18446 (n_8837, n9866);
  and g18447 (n9868, n_8836, n_8837);
  not g18448 (n_8838, n9867);
  not g18449 (n_8839, n9868);
  and g18450 (n9869, n_8838, n_8839);
  and g18451 (n9870, n_8802, n_8803);
  not g18452 (n_8840, n9870);
  and g18453 (n9871, n_8799, n_8840);
  and g18454 (n9872, n9654, n9809);
  not g18455 (n_8841, n9654);
  not g18456 (n_8842, n9809);
  and g18457 (n9873, n_8841, n_8842);
  not g18458 (n_8843, n9872);
  not g18459 (n_8844, n9873);
  and g18460 (n9874, n_8843, n_8844);
  not g18461 (n_8845, n9874);
  and g18462 (n9875, n9625, n_8845);
  not g18463 (n_8846, n9625);
  and g18464 (n9876, n_8846, n9874);
  not g18465 (n_8847, n9875);
  not g18466 (n_8848, n9876);
  and g18467 (n9877, n_8847, n_8848);
  and g18468 (n9878, n9712, n9727);
  not g18469 (n_8849, n9712);
  not g18470 (n_8850, n9727);
  and g18471 (n9879, n_8849, n_8850);
  not g18472 (n_8851, n9878);
  not g18473 (n_8852, n9879);
  and g18474 (n9880, n_8851, n_8852);
  not g18475 (n_8853, n9880);
  and g18476 (n9881, n9671, n_8853);
  not g18477 (n_8854, n9671);
  and g18478 (n9882, n_8854, n9880);
  not g18479 (n_8855, n9881);
  not g18480 (n_8856, n9882);
  and g18481 (n9883, n_8855, n_8856);
  not g18482 (n_8857, n9877);
  not g18483 (n_8858, n9883);
  and g18484 (n9884, n_8857, n_8858);
  and g18485 (n9885, n9877, n9883);
  not g18486 (n_8859, n9884);
  not g18487 (n_8860, n9885);
  and g18488 (n9886, n_8859, n_8860);
  not g18489 (n_8861, n9871);
  and g18490 (n9887, n_8861, n9886);
  not g18491 (n_8862, n9886);
  and g18492 (n9888, n9871, n_8862);
  not g18493 (n_8863, n9887);
  not g18494 (n_8864, n9888);
  and g18495 (n9889, n_8863, n_8864);
  not g18496 (n_8865, n9869);
  not g18497 (n_8866, n9889);
  and g18498 (n9890, n_8865, n_8866);
  and g18499 (n9891, n9869, n9889);
  not g18500 (n_8867, n9890);
  not g18501 (n_8868, n9891);
  and g18502 (n9892, n_8867, n_8868);
  not g18503 (n_8869, n9863);
  and g18504 (n9893, n_8869, n9892);
  not g18505 (n_8870, n9892);
  and g18506 (n9894, n9863, n_8870);
  not g18507 (n_8871, n9893);
  not g18508 (n_8872, n9894);
  and g18509 (n9895, n_8871, n_8872);
  not g18510 (n_8873, n9862);
  and g18511 (n9896, n_8873, n9895);
  not g18512 (n_8874, n9895);
  and g18513 (n9897, n9862, n_8874);
  not g18514 (n_8875, n9896);
  not g18515 (n_8876, n9897);
  and g18516 (n9898, n_8875, n_8876);
  not g18517 (n_8877, n9898);
  and g18518 (n9899, n9861, n_8877);
  not g18519 (n_8878, n9861);
  and g18520 (n9900, n_8878, n9898);
  not g18521 (n_8879, n9899);
  not g18522 (n_8880, n9900);
  and g18523 (n9901, n_8879, n_8880);
  and g18524 (n9902, n_8600, n_8605);
  and g18525 (n9903, n_8727, n_8731);
  and g18526 (n9904, n_8694, n_8695);
  not g18527 (n_8881, n9904);
  and g18528 (n9905, n_8710, n_8881);
  and g18529 (n9906, n9903, n9905);
  not g18530 (n_8882, n9903);
  not g18531 (n_8883, n9905);
  and g18532 (n9907, n_8882, n_8883);
  not g18533 (n_8884, n9906);
  not g18534 (n_8885, n9907);
  and g18535 (n9908, n_8884, n_8885);
  and g18536 (n9909, \a[61] , \a[63] );
  and g18537 (n9910, n252, n9909);
  not g18538 (n_8886, n9910);
  and g18539 (n9911, \a[61] , n_8886);
  and g18540 (n9912, \a[4] , n9911);
  and g18541 (n9913, \a[2] , n_8886);
  and g18542 (n9914, \a[63] , n9913);
  not g18543 (n_8887, n9912);
  not g18544 (n_8888, n9914);
  and g18545 (n9915, n_8887, n_8888);
  not g18546 (n_8889, n9698);
  not g18547 (n_8890, n9915);
  and g18548 (n9916, n_8889, n_8890);
  not g18549 (n_8891, n9916);
  and g18550 (n9917, n_8889, n_8891);
  and g18551 (n9918, n_8890, n_8891);
  not g18552 (n_8892, n9917);
  not g18553 (n_8893, n9918);
  and g18554 (n9919, n_8892, n_8893);
  and g18555 (n9920, n748, n7433);
  and g18556 (n9921, n8160, n8564);
  not g18557 (n_8894, n9920);
  not g18558 (n_8895, n9921);
  and g18559 (n9922, n_8894, n_8895);
  and g18560 (n9923, \a[13] , \a[52] );
  and g18561 (n9924, \a[18] , \a[47] );
  and g18562 (n9925, n9923, n9924);
  not g18563 (n_8896, n9922);
  not g18564 (n_8897, n9925);
  and g18565 (n9926, n_8896, n_8897);
  not g18566 (n_8898, n9926);
  and g18567 (n9927, n_8897, n_8898);
  not g18568 (n_8899, n9923);
  not g18569 (n_8900, n9924);
  and g18570 (n9928, n_8899, n_8900);
  not g18571 (n_8901, n9928);
  and g18572 (n9929, n9927, n_8901);
  and g18573 (n9930, \a[53] , n_8898);
  and g18574 (n9931, \a[12] , n9930);
  not g18575 (n_8902, n9929);
  not g18576 (n_8903, n9931);
  and g18577 (n9932, n_8902, n_8903);
  and g18578 (n9933, n895, n6564);
  and g18579 (n9934, \a[49] , \a[51] );
  and g18580 (n9935, n893, n9934);
  and g18581 (n9936, n891, n6325);
  not g18582 (n_8904, n9935);
  not g18583 (n_8905, n9936);
  and g18584 (n9937, n_8904, n_8905);
  not g18585 (n_8906, n9933);
  not g18586 (n_8907, n9937);
  and g18587 (n9938, n_8906, n_8907);
  not g18588 (n_8908, n9938);
  and g18589 (n9939, n7639, n_8908);
  and g18590 (n9940, \a[14] , \a[51] );
  and g18591 (n9941, \a[15] , \a[50] );
  not g18592 (n_8909, n9940);
  not g18593 (n_8910, n9941);
  and g18594 (n9942, n_8909, n_8910);
  and g18595 (n9943, n_8906, n_8908);
  not g18596 (n_8911, n9942);
  and g18597 (n9944, n_8911, n9943);
  not g18598 (n_8912, n9939);
  not g18599 (n_8913, n9944);
  and g18600 (n9945, n_8912, n_8913);
  not g18601 (n_8914, n9932);
  not g18602 (n_8915, n9945);
  and g18603 (n9946, n_8914, n_8915);
  not g18604 (n_8916, n9946);
  and g18605 (n9947, n_8914, n_8916);
  and g18606 (n9948, n_8915, n_8916);
  not g18607 (n_8917, n9947);
  not g18608 (n_8918, n9948);
  and g18609 (n9949, n_8917, n_8918);
  not g18610 (n_8919, n9919);
  and g18611 (n9950, n_8919, n9949);
  not g18612 (n_8920, n9949);
  and g18613 (n9951, n9919, n_8920);
  not g18614 (n_8921, n9950);
  not g18615 (n_8922, n9951);
  and g18616 (n9952, n_8921, n_8922);
  not g18617 (n_8923, n9952);
  and g18618 (n9953, n9908, n_8923);
  not g18619 (n_8924, n9953);
  and g18620 (n9954, n9908, n_8924);
  and g18621 (n9955, n_8923, n_8924);
  not g18622 (n_8925, n9954);
  not g18623 (n_8926, n9955);
  and g18624 (n9956, n_8925, n_8926);
  and g18625 (n9957, n9637, n9682);
  not g18626 (n_8927, n9637);
  not g18627 (n_8928, n9682);
  and g18628 (n9958, n_8927, n_8928);
  not g18629 (n_8929, n9957);
  not g18630 (n_8930, n9958);
  and g18631 (n9959, n_8929, n_8930);
  not g18632 (n_8931, n9959);
  and g18633 (n9960, n9825, n_8931);
  not g18634 (n_8932, n9825);
  and g18635 (n9961, n_8932, n9959);
  not g18636 (n_8933, n9960);
  not g18637 (n_8934, n9961);
  and g18638 (n9962, n_8933, n_8934);
  and g18639 (n9963, n_8672, n_8684);
  not g18640 (n_8935, n9962);
  and g18641 (n9964, n_8935, n9963);
  not g18642 (n_8936, n9963);
  and g18643 (n9965, n9962, n_8936);
  not g18644 (n_8937, n9964);
  not g18645 (n_8938, n9965);
  and g18646 (n9966, n_8937, n_8938);
  and g18647 (n9967, n_8635, n_8650);
  not g18648 (n_8939, n9966);
  and g18649 (n9968, n_8939, n9967);
  not g18650 (n_8940, n9967);
  and g18651 (n9969, n9966, n_8940);
  not g18652 (n_8941, n9968);
  not g18653 (n_8942, n9969);
  and g18654 (n9970, n_8941, n_8942);
  and g18655 (n9971, n_8734, n_8740);
  not g18656 (n_8943, n9971);
  and g18657 (n9972, n9970, n_8943);
  not g18658 (n_8944, n9972);
  and g18659 (n9973, n9970, n_8944);
  and g18660 (n9974, n_8943, n_8944);
  not g18661 (n_8945, n9973);
  not g18662 (n_8946, n9974);
  and g18663 (n9975, n_8945, n_8946);
  not g18664 (n_8947, n9956);
  not g18665 (n_8948, n9975);
  and g18666 (n9976, n_8947, n_8948);
  not g18667 (n_8949, n9976);
  and g18668 (n9977, n_8947, n_8949);
  and g18669 (n9978, n_8948, n_8949);
  not g18670 (n_8950, n9977);
  not g18671 (n_8951, n9978);
  and g18672 (n9979, n_8950, n_8951);
  not g18673 (n_8952, n9902);
  not g18674 (n_8953, n9979);
  and g18675 (n9980, n_8952, n_8953);
  not g18676 (n_8954, n9980);
  and g18677 (n9981, n_8952, n_8954);
  and g18678 (n9982, n_8953, n_8954);
  not g18679 (n_8955, n9981);
  not g18680 (n_8956, n9982);
  and g18681 (n9983, n_8955, n_8956);
  and g18682 (n9984, n_8569, n_8598);
  and g18683 (n9985, \a[20] , \a[56] );
  and g18684 (n9986, n6997, n9985);
  and g18685 (n9987, n484, n9161);
  not g18686 (n_8957, n9986);
  not g18687 (n_8958, n9987);
  and g18688 (n9988, n_8957, n_8958);
  and g18689 (n9989, \a[10] , \a[55] );
  and g18690 (n9990, \a[20] , \a[45] );
  and g18691 (n9991, n9989, n9990);
  not g18692 (n_8959, n9988);
  not g18693 (n_8960, n9991);
  and g18694 (n9992, n_8959, n_8960);
  not g18695 (n_8961, n9992);
  and g18696 (n9993, n_8960, n_8961);
  not g18697 (n_8962, n9989);
  not g18698 (n_8963, n9990);
  and g18699 (n9994, n_8962, n_8963);
  not g18700 (n_8964, n9994);
  and g18701 (n9995, n9993, n_8964);
  and g18702 (n9996, \a[56] , n_8961);
  and g18703 (n9997, \a[9] , n9996);
  not g18704 (n_8965, n9995);
  not g18705 (n_8966, n9997);
  and g18706 (n9998, n_8965, n_8966);
  and g18707 (n9999, n1904, n5413);
  and g18708 (n10000, n1547, n6453);
  and g18709 (n10001, n1666, n5344);
  not g18710 (n_8967, n10000);
  not g18711 (n_8968, n10001);
  and g18712 (n10002, n_8967, n_8968);
  not g18713 (n_8969, n9999);
  not g18714 (n_8970, n10002);
  and g18715 (n10003, n_8969, n_8970);
  not g18716 (n_8971, n10003);
  and g18717 (n10004, \a[42] , n_8971);
  and g18718 (n10005, \a[23] , n10004);
  and g18719 (n10006, \a[24] , \a[41] );
  and g18720 (n10007, \a[25] , \a[40] );
  not g18721 (n_8972, n10006);
  not g18722 (n_8973, n10007);
  and g18723 (n10008, n_8972, n_8973);
  and g18724 (n10009, n_8969, n_8971);
  not g18725 (n_8974, n10008);
  and g18726 (n10010, n_8974, n10009);
  not g18727 (n_8975, n10005);
  not g18728 (n_8976, n10010);
  and g18729 (n10011, n_8975, n_8976);
  not g18730 (n_8977, n9998);
  not g18731 (n_8978, n10011);
  and g18732 (n10012, n_8977, n_8978);
  not g18733 (n_8979, n10012);
  and g18734 (n10013, n_8977, n_8979);
  and g18735 (n10014, n_8978, n_8979);
  not g18736 (n_8980, n10013);
  not g18737 (n_8981, n10014);
  and g18738 (n10015, n_8980, n_8981);
  and g18739 (n10016, n2331, n4565);
  and g18740 (n10017, n2800, n5430);
  and g18741 (n10018, n2227, n5083);
  not g18742 (n_8982, n10017);
  not g18743 (n_8983, n10018);
  and g18744 (n10019, n_8982, n_8983);
  not g18745 (n_8984, n10016);
  not g18746 (n_8985, n10019);
  and g18747 (n10020, n_8984, n_8985);
  not g18748 (n_8986, n10020);
  and g18749 (n10021, \a[39] , n_8986);
  and g18750 (n10022, \a[26] , n10021);
  and g18751 (n10023, n_8984, n_8986);
  and g18752 (n10024, \a[27] , \a[38] );
  and g18753 (n10025, \a[28] , \a[37] );
  not g18754 (n_8987, n10024);
  not g18755 (n_8988, n10025);
  and g18756 (n10026, n_8987, n_8988);
  not g18757 (n_8989, n10026);
  and g18758 (n10027, n10023, n_8989);
  not g18759 (n_8990, n10022);
  not g18760 (n_8991, n10027);
  and g18761 (n10028, n_8990, n_8991);
  not g18762 (n_8992, n10015);
  not g18763 (n_8993, n10028);
  and g18764 (n10029, n_8992, n_8993);
  not g18765 (n_8994, n10029);
  and g18766 (n10030, n_8992, n_8994);
  and g18767 (n10031, n_8993, n_8994);
  not g18768 (n_8995, n10030);
  not g18769 (n_8996, n10031);
  and g18770 (n10032, n_8995, n_8996);
  and g18771 (n10033, \a[11] , \a[54] );
  and g18772 (n10034, \a[19] , \a[46] );
  not g18773 (n_8997, n10033);
  not g18774 (n_8998, n10034);
  and g18775 (n10035, n_8997, n_8998);
  and g18776 (n10036, n10033, n10034);
  not g18777 (n_8999, n10036);
  not g18780 (n_9000, n10035);
  not g18782 (n_9001, n10039);
  and g18783 (n10040, n_8999, n_9001);
  and g18784 (n10041, n_9000, n10040);
  and g18785 (n10042, \a[36] , n_9001);
  and g18786 (n10043, \a[29] , n10042);
  not g18787 (n_9002, n10041);
  not g18788 (n_9003, n10043);
  and g18789 (n10044, n_9002, n_9003);
  and g18790 (n10045, n3812, n4150);
  and g18791 (n10046, n3143, n4024);
  and g18792 (n10047, n2865, n3319);
  not g18793 (n_9004, n10046);
  not g18794 (n_9005, n10047);
  and g18795 (n10048, n_9004, n_9005);
  not g18796 (n_9006, n10045);
  not g18797 (n_9007, n10048);
  and g18798 (n10049, n_9006, n_9007);
  not g18799 (n_9008, n10049);
  and g18800 (n10050, n4024, n_9008);
  and g18801 (n10051, n_9006, n_9008);
  not g18802 (n_9009, n3143);
  not g18803 (n_9010, n6485);
  and g18804 (n10052, n_9009, n_9010);
  not g18805 (n_9011, n10052);
  and g18806 (n10053, n10051, n_9011);
  not g18807 (n_9012, n10050);
  not g18808 (n_9013, n10053);
  and g18809 (n10054, n_9012, n_9013);
  not g18810 (n_9014, n10044);
  not g18811 (n_9015, n10054);
  and g18812 (n10055, n_9014, n_9015);
  not g18813 (n_9016, n10055);
  and g18814 (n10056, n_9014, n_9016);
  and g18815 (n10057, n_9015, n_9016);
  not g18816 (n_9017, n10056);
  not g18817 (n_9018, n10057);
  and g18818 (n10058, n_9017, n_9018);
  and g18819 (n10059, \a[3] , \a[62] );
  not g18820 (n_9019, \a[33] );
  not g18821 (n_9020, n10059);
  and g18822 (n10060, n_9019, n_9020);
  and g18823 (n10061, \a[33] , n10059);
  not g18824 (n_9021, n10061);
  and g18825 (n10062, n6944, n_9021);
  not g18826 (n_9022, n10060);
  and g18827 (n10063, n_9022, n10062);
  not g18828 (n_9023, n10063);
  and g18829 (n10064, n6944, n_9023);
  and g18830 (n10065, n_9021, n_9023);
  and g18831 (n10066, n_9022, n10065);
  not g18832 (n_9024, n10064);
  not g18833 (n_9025, n10066);
  and g18834 (n10067, n_9024, n_9025);
  not g18835 (n_9026, n10058);
  not g18836 (n_9027, n10067);
  and g18837 (n10068, n_9026, n_9027);
  not g18838 (n_9028, n10068);
  and g18839 (n10069, n_9026, n_9028);
  and g18840 (n10070, n_9027, n_9028);
  not g18841 (n_9029, n10069);
  not g18842 (n_9030, n10070);
  and g18843 (n10071, n_9029, n_9030);
  and g18844 (n10072, \a[21] , \a[44] );
  and g18845 (n10073, \a[22] , \a[43] );
  not g18846 (n_9031, n10072);
  not g18847 (n_9032, n10073);
  and g18848 (n10074, n_9031, n_9032);
  and g18849 (n10075, n1574, n5296);
  not g18850 (n_9033, n10075);
  not g18853 (n_9034, n10074);
  not g18855 (n_9035, n10078);
  and g18856 (n10079, \a[8] , n_9035);
  and g18857 (n10080, \a[57] , n10079);
  and g18858 (n10081, n_9033, n_9035);
  and g18859 (n10082, n_9034, n10081);
  not g18860 (n_9036, n10080);
  not g18861 (n_9037, n10082);
  and g18862 (n10083, n_9036, n_9037);
  and g18863 (n10084, n_8769, n_8774);
  not g18864 (n_9038, n10083);
  and g18865 (n10085, n_9038, n10084);
  not g18866 (n_9039, n10084);
  and g18867 (n10086, n10083, n_9039);
  not g18868 (n_9040, n10085);
  not g18869 (n_9041, n10086);
  and g18870 (n10087, n_9040, n_9041);
  and g18871 (n10088, n335, n8987);
  and g18872 (n10089, \a[58] , \a[60] );
  and g18873 (n10090, n268, n10089);
  and g18874 (n10091, n332, n9509);
  not g18875 (n_9042, n10090);
  not g18876 (n_9043, n10091);
  and g18877 (n10092, n_9042, n_9043);
  not g18878 (n_9044, n10088);
  not g18879 (n_9045, n10092);
  and g18880 (n10093, n_9044, n_9045);
  not g18881 (n_9046, n10093);
  and g18882 (n10094, \a[60] , n_9046);
  and g18883 (n10095, \a[5] , n10094);
  and g18884 (n10096, n_9044, n_9046);
  and g18885 (n10097, \a[6] , \a[59] );
  and g18886 (n10098, \a[7] , \a[58] );
  not g18887 (n_9047, n10097);
  not g18888 (n_9048, n10098);
  and g18889 (n10099, n_9047, n_9048);
  not g18890 (n_9049, n10099);
  and g18891 (n10100, n10096, n_9049);
  not g18892 (n_9050, n10095);
  not g18893 (n_9051, n10100);
  and g18894 (n10101, n_9050, n_9051);
  not g18895 (n_9052, n10087);
  not g18896 (n_9053, n10101);
  and g18897 (n10102, n_9052, n_9053);
  and g18898 (n10103, n10087, n10101);
  not g18899 (n_9054, n10102);
  not g18900 (n_9055, n10103);
  and g18901 (n10104, n_9054, n_9055);
  and g18902 (n10105, n10071, n10104);
  not g18903 (n_9056, n10071);
  not g18904 (n_9057, n10104);
  and g18905 (n10106, n_9056, n_9057);
  not g18906 (n_9058, n10105);
  not g18907 (n_9059, n10106);
  and g18908 (n10107, n_9058, n_9059);
  not g18909 (n_9060, n10032);
  not g18910 (n_9061, n10107);
  and g18911 (n10108, n_9060, n_9061);
  not g18912 (n_9062, n10108);
  and g18913 (n10109, n_9060, n_9062);
  and g18914 (n10110, n_9061, n_9062);
  not g18915 (n_9063, n10109);
  not g18916 (n_9064, n10110);
  and g18917 (n10111, n_9063, n_9064);
  not g18918 (n_9065, n9984);
  not g18919 (n_9066, n10111);
  and g18920 (n10112, n_9065, n_9066);
  not g18921 (n_9067, n10112);
  and g18922 (n10113, n_9065, n_9067);
  and g18923 (n10114, n_9066, n_9067);
  not g18924 (n_9068, n10113);
  not g18925 (n_9069, n10114);
  and g18926 (n10115, n_9068, n_9069);
  and g18927 (n10116, n_8747, n_8751);
  and g18928 (n10117, n_8574, n_8578);
  and g18929 (n10118, n10116, n10117);
  not g18930 (n_9070, n10116);
  not g18931 (n_9071, n10117);
  and g18932 (n10119, n_9070, n_9071);
  not g18933 (n_9072, n10118);
  not g18934 (n_9073, n10119);
  and g18935 (n10120, n_9072, n_9073);
  and g18936 (n10121, n_8582, n_8586);
  not g18937 (n_9074, n10120);
  and g18938 (n10122, n_9074, n10121);
  not g18939 (n_9075, n10121);
  and g18940 (n10123, n10120, n_9075);
  not g18941 (n_9076, n10122);
  not g18942 (n_9077, n10123);
  and g18943 (n10124, n_9076, n_9077);
  and g18944 (n10125, n_8590, n_8593);
  and g18945 (n10126, n_8755, n_8759);
  not g18946 (n_9078, n10125);
  and g18947 (n10127, n_9078, n10126);
  not g18948 (n_9079, n10126);
  and g18949 (n10128, n10125, n_9079);
  not g18950 (n_9080, n10127);
  not g18951 (n_9081, n10128);
  and g18952 (n10129, n_9080, n_9081);
  not g18953 (n_9082, n10129);
  and g18954 (n10130, n10124, n_9082);
  not g18955 (n_9083, n10124);
  and g18956 (n10131, n_9083, n10129);
  not g18957 (n_9084, n10130);
  not g18958 (n_9085, n10131);
  and g18959 (n10132, n_9084, n_9085);
  not g18960 (n_9086, n10115);
  and g18961 (n10133, n_9086, n10132);
  not g18962 (n_9087, n10133);
  and g18963 (n10134, n_9086, n_9087);
  and g18964 (n10135, n10132, n_9087);
  not g18965 (n_9088, n10134);
  not g18966 (n_9089, n10135);
  and g18967 (n10136, n_9088, n_9089);
  not g18968 (n_9090, n9983);
  and g18969 (n10137, n_9090, n10136);
  not g18970 (n_9091, n10136);
  and g18971 (n10138, n9983, n_9091);
  not g18972 (n_9092, n10137);
  not g18973 (n_9093, n10138);
  and g18974 (n10139, n_9092, n_9093);
  not g18975 (n_9094, n10139);
  and g18976 (n10140, n9901, n_9094);
  not g18977 (n_9095, n9901);
  and g18978 (n10141, n_9095, n10139);
  not g18979 (n_9096, n10140);
  not g18980 (n_9097, n10141);
  and g18981 (n10142, n_9096, n_9097);
  not g18982 (n_9098, n9860);
  and g18983 (n10143, n_9098, n10142);
  not g18984 (n_9099, n10142);
  and g18985 (n10144, n9860, n_9099);
  not g18986 (n_9100, n10143);
  not g18987 (n_9101, n10144);
  and g18988 (n10145, n_9100, n_9101);
  not g18989 (n_9102, n9859);
  not g18990 (n_9103, n10145);
  and g18991 (n10146, n_9102, n_9103);
  and g18992 (n10147, n9859, n10145);
  or g18993 (\asquared[66] , n10146, n10147);
  and g18994 (n10149, n_9102, n_9101);
  not g18995 (n_9104, n10149);
  and g18996 (n10150, n_9100, n_9104);
  and g18997 (n10151, n_8880, n_9096);
  and g18998 (n10152, n_9090, n_9091);
  not g18999 (n_9105, n10152);
  and g19000 (n10153, n_8954, n_9105);
  and g19001 (n10154, n_8944, n_8949);
  and g19002 (n10155, n9927, n9993);
  not g19003 (n_9106, n9927);
  not g19004 (n_9107, n9993);
  and g19005 (n10156, n_9106, n_9107);
  not g19006 (n_9108, n10155);
  not g19007 (n_9109, n10156);
  and g19008 (n10157, n_9108, n_9109);
  not g19009 (n_9110, n10157);
  and g19010 (n10158, n10009, n_9110);
  not g19011 (n_9111, n10009);
  and g19012 (n10159, n_9111, n10157);
  not g19013 (n_9112, n10158);
  not g19014 (n_9113, n10159);
  and g19015 (n10160, n_9112, n_9113);
  and g19016 (n10161, n_9038, n_9039);
  not g19017 (n_9114, n10161);
  and g19018 (n10162, n_9054, n_9114);
  not g19019 (n_9115, n10160);
  and g19020 (n10163, n_9115, n10162);
  not g19021 (n_9116, n10162);
  and g19022 (n10164, n10160, n_9116);
  not g19023 (n_9117, n10163);
  not g19024 (n_9118, n10164);
  and g19025 (n10165, n_9117, n_9118);
  and g19026 (n10166, n_8979, n_8994);
  not g19027 (n_9119, n10165);
  and g19028 (n10167, n_9119, n10166);
  not g19029 (n_9120, n10166);
  and g19030 (n10168, n10165, n_9120);
  not g19031 (n_9121, n10167);
  not g19032 (n_9122, n10168);
  and g19033 (n10169, n_9121, n_9122);
  and g19034 (n10170, n_9056, n10104);
  not g19035 (n_9123, n10170);
  and g19036 (n10171, n_9062, n_9123);
  and g19037 (n10172, n_8885, n_8924);
  and g19038 (n10173, n10171, n10172);
  not g19039 (n_9124, n10171);
  not g19040 (n_9125, n10172);
  and g19041 (n10174, n_9124, n_9125);
  not g19042 (n_9126, n10173);
  not g19043 (n_9127, n10174);
  and g19044 (n10175, n_9126, n_9127);
  and g19045 (n10176, n10169, n10175);
  not g19046 (n_9128, n10169);
  not g19047 (n_9129, n10175);
  and g19048 (n10177, n_9128, n_9129);
  not g19049 (n_9130, n10176);
  not g19050 (n_9131, n10177);
  and g19051 (n10178, n_9130, n_9131);
  not g19052 (n_9132, n10154);
  and g19053 (n10179, n_9132, n10178);
  not g19054 (n_9133, n10179);
  and g19055 (n10180, n_9132, n_9133);
  and g19056 (n10181, n10178, n_9133);
  not g19057 (n_9134, n10180);
  not g19058 (n_9135, n10181);
  and g19059 (n10182, n_9134, n_9135);
  and g19060 (n10183, n_9078, n_9079);
  not g19061 (n_9136, n10183);
  and g19062 (n10184, n_9084, n_9136);
  and g19063 (n10185, n_8886, n_8891);
  and g19064 (n10186, n10023, n10185);
  not g19065 (n_9137, n10023);
  not g19066 (n_9138, n10185);
  and g19067 (n10187, n_9137, n_9138);
  not g19068 (n_9139, n10186);
  not g19069 (n_9140, n10187);
  and g19070 (n10188, n_9139, n_9140);
  and g19071 (n10189, n380, n8987);
  and g19072 (n10190, n312, n10089);
  and g19073 (n10191, n335, n9509);
  not g19074 (n_9141, n10190);
  not g19075 (n_9142, n10191);
  and g19076 (n10192, n_9141, n_9142);
  not g19077 (n_9143, n10189);
  not g19078 (n_9144, n10192);
  and g19079 (n10193, n_9143, n_9144);
  not g19080 (n_9145, n10193);
  and g19081 (n10194, \a[60] , n_9145);
  and g19082 (n10195, \a[6] , n10194);
  and g19083 (n10196, n_9143, n_9145);
  and g19084 (n10197, \a[7] , \a[59] );
  and g19085 (n10198, \a[8] , \a[58] );
  not g19086 (n_9146, n10197);
  not g19087 (n_9147, n10198);
  and g19088 (n10199, n_9146, n_9147);
  not g19089 (n_9148, n10199);
  and g19090 (n10200, n10196, n_9148);
  not g19091 (n_9149, n10195);
  not g19092 (n_9150, n10200);
  and g19093 (n10201, n_9149, n_9150);
  not g19094 (n_9151, n10201);
  and g19095 (n10202, n10188, n_9151);
  not g19096 (n_9152, n10202);
  and g19097 (n10203, n10188, n_9152);
  and g19098 (n10204, n_9151, n_9152);
  not g19099 (n_9153, n10203);
  not g19100 (n_9154, n10204);
  and g19101 (n10205, n_9153, n_9154);
  and g19102 (n10206, n_8919, n_8920);
  not g19103 (n_9155, n10206);
  and g19104 (n10207, n_8916, n_9155);
  not g19105 (n_9156, n10205);
  not g19106 (n_9157, n10207);
  and g19107 (n10208, n_9156, n_9157);
  not g19108 (n_9158, n10208);
  and g19109 (n10209, n_9156, n_9158);
  and g19110 (n10210, n_9157, n_9158);
  not g19111 (n_9159, n10209);
  not g19112 (n_9160, n10210);
  and g19113 (n10211, n_9159, n_9160);
  and g19114 (n10212, n_9073, n_9077);
  and g19115 (n10213, n10211, n10212);
  not g19116 (n_9161, n10211);
  not g19117 (n_9162, n10212);
  and g19118 (n10214, n_9161, n_9162);
  not g19119 (n_9163, n10213);
  not g19120 (n_9164, n10214);
  and g19121 (n10215, n_9163, n_9164);
  and g19122 (n10216, n10051, n10065);
  not g19123 (n_9165, n10051);
  not g19124 (n_9166, n10065);
  and g19125 (n10217, n_9165, n_9166);
  not g19126 (n_9167, n10216);
  not g19127 (n_9168, n10217);
  and g19128 (n10218, n_9167, n_9168);
  not g19129 (n_9169, n10218);
  and g19130 (n10219, n9943, n_9169);
  not g19131 (n_9170, n9943);
  and g19132 (n10220, n_9170, n10218);
  not g19133 (n_9171, n10219);
  not g19134 (n_9172, n10220);
  and g19135 (n10221, n_9171, n_9172);
  and g19136 (n10222, n10081, n10096);
  not g19137 (n_9173, n10081);
  not g19138 (n_9174, n10096);
  and g19139 (n10223, n_9173, n_9174);
  not g19140 (n_9175, n10222);
  not g19141 (n_9176, n10223);
  and g19142 (n10224, n_9175, n_9176);
  not g19143 (n_9177, n10224);
  and g19144 (n10225, n10040, n_9177);
  not g19145 (n_9178, n10040);
  and g19146 (n10226, n_9178, n10224);
  not g19147 (n_9179, n10225);
  not g19148 (n_9180, n10226);
  and g19149 (n10227, n_9179, n_9180);
  and g19150 (n10228, n_9016, n_9028);
  not g19151 (n_9181, n10227);
  and g19152 (n10229, n_9181, n10228);
  not g19153 (n_9182, n10228);
  and g19154 (n10230, n10227, n_9182);
  not g19155 (n_9183, n10229);
  not g19156 (n_9184, n10230);
  and g19157 (n10231, n_9183, n_9184);
  and g19158 (n10232, n10221, n10231);
  not g19159 (n_9185, n10221);
  not g19160 (n_9186, n10231);
  and g19161 (n10233, n_9185, n_9186);
  not g19162 (n_9187, n10232);
  not g19163 (n_9188, n10233);
  and g19164 (n10234, n_9187, n_9188);
  and g19165 (n10235, n10215, n10234);
  not g19166 (n_9189, n10215);
  not g19167 (n_9190, n10234);
  and g19168 (n10236, n_9189, n_9190);
  not g19169 (n_9191, n10235);
  not g19170 (n_9192, n10236);
  and g19171 (n10237, n_9191, n_9192);
  not g19172 (n_9193, n10184);
  and g19173 (n10238, n_9193, n10237);
  not g19174 (n_9194, n10237);
  and g19175 (n10239, n10184, n_9194);
  not g19176 (n_9195, n10238);
  not g19177 (n_9196, n10239);
  and g19178 (n10240, n_9195, n_9196);
  not g19179 (n_9197, n10182);
  and g19180 (n10241, n_9197, n10240);
  not g19181 (n_9198, n10241);
  and g19182 (n10242, n10240, n_9198);
  and g19183 (n10243, n_9197, n_9198);
  not g19184 (n_9199, n10242);
  not g19185 (n_9200, n10243);
  and g19186 (n10244, n_9199, n_9200);
  not g19187 (n_9201, n10153);
  not g19188 (n_9202, n10244);
  and g19189 (n10245, n_9201, n_9202);
  not g19190 (n_9203, n10245);
  and g19191 (n10246, n_9201, n_9203);
  and g19192 (n10247, n_9202, n_9203);
  not g19193 (n_9204, n10246);
  not g19194 (n_9205, n10247);
  and g19195 (n10248, n_9204, n_9205);
  and g19196 (n10249, n_8871, n_8875);
  and g19197 (n10250, n_9067, n_9087);
  and g19198 (n10251, n10249, n10250);
  not g19199 (n_9206, n10249);
  not g19200 (n_9207, n10250);
  and g19201 (n10252, n_9206, n_9207);
  not g19202 (n_9208, n10251);
  not g19203 (n_9209, n10252);
  and g19204 (n10253, n_9208, n_9209);
  and g19205 (n10254, n_8839, n_8868);
  and g19206 (n10255, n226, n9721);
  and g19207 (n10256, n300, n9909);
  and g19208 (n10257, n209, n9792);
  not g19209 (n_9210, n10256);
  not g19210 (n_9211, n10257);
  and g19211 (n10258, n_9210, n_9211);
  not g19212 (n_9212, n10255);
  not g19213 (n_9213, n10258);
  and g19214 (n10259, n_9212, n_9213);
  not g19215 (n_9214, n10259);
  and g19216 (n10260, n_9212, n_9214);
  and g19217 (n10261, \a[4] , \a[62] );
  not g19218 (n_9215, n8907);
  not g19219 (n_9216, n10261);
  and g19220 (n10262, n_9215, n_9216);
  not g19221 (n_9217, n10262);
  and g19222 (n10263, n10260, n_9217);
  and g19223 (n10264, \a[63] , n_9214);
  and g19224 (n10265, \a[3] , n10264);
  not g19225 (n_9218, n10263);
  not g19226 (n_9219, n10265);
  and g19227 (n10266, n_9218, n_9219);
  and g19228 (n10267, n2334, n4565);
  and g19229 (n10268, n2041, n5430);
  and g19230 (n10269, n2331, n5083);
  not g19231 (n_9220, n10268);
  not g19232 (n_9221, n10269);
  and g19233 (n10270, n_9220, n_9221);
  not g19234 (n_9222, n10267);
  not g19235 (n_9223, n10270);
  and g19236 (n10271, n_9222, n_9223);
  not g19237 (n_9224, n10271);
  and g19238 (n10272, \a[39] , n_9224);
  and g19239 (n10273, \a[27] , n10272);
  and g19240 (n10274, \a[28] , \a[38] );
  and g19241 (n10275, \a[29] , \a[37] );
  not g19242 (n_9225, n10274);
  not g19243 (n_9226, n10275);
  and g19244 (n10276, n_9225, n_9226);
  and g19245 (n10277, n_9222, n_9224);
  not g19246 (n_9227, n10276);
  and g19247 (n10278, n_9227, n10277);
  not g19248 (n_9228, n10273);
  not g19249 (n_9229, n10278);
  and g19250 (n10279, n_9228, n_9229);
  not g19251 (n_9230, n10266);
  not g19252 (n_9231, n10279);
  and g19253 (n10280, n_9230, n_9231);
  not g19254 (n_9232, n10280);
  and g19255 (n10281, n_9230, n_9232);
  and g19256 (n10282, n_9231, n_9232);
  not g19257 (n_9233, n10281);
  not g19258 (n_9234, n10282);
  and g19259 (n10283, n_9233, n_9234);
  and g19260 (n10284, \a[19] , \a[47] );
  and g19261 (n10285, \a[12] , \a[54] );
  and g19262 (n10286, n10284, n10285);
  and g19263 (n10287, n602, n7701);
  and g19264 (n10288, n8060, n8212);
  not g19265 (n_9235, n10287);
  not g19266 (n_9236, n10288);
  and g19267 (n10289, n_9235, n_9236);
  not g19268 (n_9237, n10286);
  not g19269 (n_9238, n10289);
  and g19270 (n10290, n_9237, n_9238);
  not g19271 (n_9239, n10290);
  and g19272 (n10291, \a[55] , n_9239);
  and g19273 (n10292, \a[11] , n10291);
  and g19274 (n10293, n_9237, n_9239);
  not g19275 (n_9240, n10284);
  not g19276 (n_9241, n10285);
  and g19277 (n10294, n_9240, n_9241);
  not g19278 (n_9242, n10294);
  and g19279 (n10295, n10293, n_9242);
  not g19280 (n_9243, n10292);
  not g19281 (n_9244, n10295);
  and g19282 (n10296, n_9243, n_9244);
  not g19283 (n_9245, n10283);
  not g19284 (n_9246, n10296);
  and g19285 (n10297, n_9245, n_9246);
  not g19286 (n_9247, n10297);
  and g19287 (n10298, n_9245, n_9247);
  and g19288 (n10299, n_9246, n_9247);
  not g19289 (n_9248, n10298);
  not g19290 (n_9249, n10299);
  and g19291 (n10300, n_9248, n_9249);
  and g19292 (n10301, \a[24] , \a[57] );
  and g19293 (n10302, n6180, n10301);
  and g19294 (n10303, \a[43] , \a[57] );
  and g19295 (n10304, \a[23] , n10303);
  and g19296 (n10305, \a[9] , n10304);
  and g19297 (n10306, n1666, n5018);
  not g19298 (n_9250, n10305);
  not g19299 (n_9251, n10306);
  and g19300 (n10307, n_9250, n_9251);
  not g19301 (n_9252, n10302);
  not g19302 (n_9253, n10307);
  and g19303 (n10308, n_9252, n_9253);
  not g19304 (n_9254, n10308);
  and g19305 (n10309, n_9252, n_9254);
  and g19306 (n10310, \a[9] , \a[57] );
  and g19307 (n10311, \a[24] , \a[42] );
  not g19308 (n_9255, n10310);
  not g19309 (n_9256, n10311);
  and g19310 (n10312, n_9255, n_9256);
  not g19311 (n_9257, n10312);
  and g19312 (n10313, n10309, n_9257);
  and g19313 (n10314, \a[43] , n_9254);
  and g19314 (n10315, \a[23] , n10314);
  not g19315 (n_9258, n10313);
  not g19316 (n_9259, n10315);
  and g19317 (n10316, n_9258, n_9259);
  and g19318 (n10317, n1574, n5713);
  and g19319 (n10318, n1693, n7747);
  and g19320 (n10319, n1494, n5560);
  not g19321 (n_9260, n10318);
  not g19322 (n_9261, n10319);
  and g19323 (n10320, n_9260, n_9261);
  not g19324 (n_9262, n10317);
  not g19325 (n_9263, n10320);
  and g19326 (n10321, n_9262, n_9263);
  not g19327 (n_9264, n10321);
  and g19328 (n10322, \a[46] , n_9264);
  and g19329 (n10323, \a[20] , n10322);
  and g19330 (n10324, \a[21] , \a[45] );
  and g19331 (n10325, \a[22] , \a[44] );
  not g19332 (n_9265, n10324);
  not g19333 (n_9266, n10325);
  and g19334 (n10326, n_9265, n_9266);
  and g19335 (n10327, n_9262, n_9264);
  not g19336 (n_9267, n10326);
  and g19337 (n10328, n_9267, n10327);
  not g19338 (n_9268, n10323);
  not g19339 (n_9269, n10328);
  and g19340 (n10329, n_9268, n_9269);
  not g19341 (n_9270, n10316);
  not g19342 (n_9271, n10329);
  and g19343 (n10330, n_9270, n_9271);
  not g19344 (n_9272, n10330);
  and g19345 (n10331, n_9270, n_9272);
  and g19346 (n10332, n_9271, n_9272);
  not g19347 (n_9273, n10331);
  not g19348 (n_9274, n10332);
  and g19349 (n10333, n_9273, n_9274);
  and g19350 (n10334, \a[25] , \a[41] );
  and g19351 (n10335, \a[26] , \a[40] );
  not g19352 (n_9275, n10334);
  not g19353 (n_9276, n10335);
  and g19354 (n10336, n_9275, n_9276);
  and g19355 (n10337, n2463, n5413);
  not g19356 (n_9277, n10337);
  not g19359 (n_9278, n10336);
  not g19361 (n_9279, n10340);
  and g19362 (n10341, \a[56] , n_9279);
  and g19363 (n10342, \a[10] , n10341);
  and g19364 (n10343, n_9277, n_9279);
  and g19365 (n10344, n_9278, n10343);
  not g19366 (n_9280, n10342);
  not g19367 (n_9281, n10344);
  and g19368 (n10345, n_9280, n_9281);
  not g19369 (n_9282, n10333);
  not g19370 (n_9283, n10345);
  and g19371 (n10346, n_9282, n_9283);
  not g19372 (n_9284, n10346);
  and g19373 (n10347, n_9282, n_9284);
  and g19374 (n10348, n_9283, n_9284);
  not g19375 (n_9285, n10347);
  not g19376 (n_9286, n10348);
  and g19377 (n10349, n_9285, n_9286);
  and g19378 (n10350, \a[13] , \a[53] );
  and g19379 (n10351, \a[15] , \a[51] );
  not g19380 (n_9287, n10350);
  not g19381 (n_9288, n10351);
  and g19382 (n10352, n_9287, n_9288);
  and g19383 (n10353, n821, n7232);
  not g19384 (n_9289, n10353);
  not g19387 (n_9290, n10352);
  not g19389 (n_9291, n10356);
  and g19390 (n10357, n_9289, n_9291);
  and g19391 (n10358, n_9290, n10357);
  and g19392 (n10359, \a[48] , n_9291);
  and g19393 (n10360, \a[18] , n10359);
  not g19394 (n_9292, n10358);
  not g19395 (n_9293, n10360);
  and g19396 (n10361, n_9292, n_9293);
  and g19397 (n10362, \a[31] , \a[35] );
  not g19398 (n_9294, n4027);
  not g19399 (n_9295, n10362);
  and g19400 (n10363, n_9294, n_9295);
  and g19401 (n10364, n2865, n3828);
  not g19402 (n_9296, n10364);
  not g19405 (n_9297, n10363);
  not g19407 (n_9298, n10367);
  and g19408 (n10368, \a[52] , n_9298);
  and g19409 (n10369, \a[14] , n10368);
  and g19410 (n10370, n_9296, n_9298);
  and g19411 (n10371, n_9297, n10370);
  not g19412 (n_9299, n10369);
  not g19413 (n_9300, n10371);
  and g19414 (n10372, n_9299, n_9300);
  not g19415 (n_9301, n10361);
  not g19416 (n_9302, n10372);
  and g19417 (n10373, n_9301, n_9302);
  not g19418 (n_9303, n10373);
  and g19419 (n10374, n_9301, n_9303);
  and g19420 (n10375, n_9302, n_9303);
  not g19421 (n_9304, n10374);
  not g19422 (n_9305, n10375);
  and g19423 (n10376, n_9304, n_9305);
  not g19424 (n_9306, n7063);
  not g19425 (n_9307, n7642);
  and g19426 (n10377, n_9306, n_9307);
  and g19427 (n10378, n1048, n6325);
  not g19428 (n_9308, n10378);
  and g19429 (n10379, n4090, n_9308);
  not g19430 (n_9309, n10377);
  and g19431 (n10380, n_9309, n10379);
  not g19432 (n_9310, n10380);
  and g19433 (n10381, n4090, n_9310);
  and g19434 (n10382, n_9308, n_9310);
  and g19435 (n10383, n_9309, n10382);
  not g19436 (n_9311, n10381);
  not g19437 (n_9312, n10383);
  and g19438 (n10384, n_9311, n_9312);
  not g19439 (n_9313, n10376);
  not g19440 (n_9314, n10384);
  and g19441 (n10385, n_9313, n_9314);
  not g19442 (n_9315, n10385);
  and g19443 (n10386, n_9313, n_9315);
  and g19444 (n10387, n_9314, n_9315);
  not g19445 (n_9316, n10386);
  not g19446 (n_9317, n10387);
  and g19447 (n10388, n_9316, n_9317);
  not g19448 (n_9318, n10349);
  and g19449 (n10389, n_9318, n10388);
  not g19450 (n_9319, n10388);
  and g19451 (n10390, n10349, n_9319);
  not g19452 (n_9320, n10389);
  not g19453 (n_9321, n10390);
  and g19454 (n10391, n_9320, n_9321);
  not g19455 (n_9322, n10300);
  not g19456 (n_9323, n10391);
  and g19457 (n10392, n_9322, n_9323);
  and g19458 (n10393, n10300, n10391);
  not g19459 (n_9324, n10392);
  not g19460 (n_9325, n10393);
  and g19461 (n10394, n_9324, n_9325);
  not g19462 (n_9326, n10254);
  and g19463 (n10395, n_9326, n10394);
  not g19464 (n_9327, n10394);
  and g19465 (n10396, n10254, n_9327);
  not g19466 (n_9328, n10395);
  not g19467 (n_9329, n10396);
  and g19468 (n10397, n_9328, n_9329);
  and g19469 (n10398, n_8844, n_8848);
  and g19470 (n10399, n_8852, n_8856);
  and g19471 (n10400, n10398, n10399);
  not g19472 (n_9330, n10398);
  not g19473 (n_9331, n10399);
  and g19474 (n10401, n_9330, n_9331);
  not g19475 (n_9332, n10400);
  not g19476 (n_9333, n10401);
  and g19477 (n10402, n_9332, n_9333);
  and g19478 (n10403, n_8930, n_8934);
  not g19479 (n_9334, n10402);
  and g19480 (n10404, n_9334, n10403);
  not g19481 (n_9335, n10403);
  and g19482 (n10405, n10402, n_9335);
  not g19483 (n_9336, n10404);
  not g19484 (n_9337, n10405);
  and g19485 (n10406, n_9336, n_9337);
  and g19486 (n10407, n_8860, n_8863);
  and g19487 (n10408, n_8938, n_8942);
  not g19488 (n_9338, n10407);
  and g19489 (n10409, n_9338, n10408);
  not g19490 (n_9339, n10408);
  and g19491 (n10410, n10407, n_9339);
  not g19492 (n_9340, n10409);
  not g19493 (n_9341, n10410);
  and g19494 (n10411, n_9340, n_9341);
  not g19495 (n_9342, n10411);
  and g19496 (n10412, n10406, n_9342);
  not g19497 (n_9343, n10406);
  and g19498 (n10413, n_9343, n10411);
  not g19499 (n_9344, n10412);
  not g19500 (n_9345, n10413);
  and g19501 (n10414, n_9344, n_9345);
  and g19502 (n10415, n10397, n10414);
  not g19503 (n_9346, n10397);
  not g19504 (n_9347, n10414);
  and g19505 (n10416, n_9346, n_9347);
  not g19506 (n_9348, n10415);
  not g19507 (n_9349, n10416);
  and g19508 (n10417, n_9348, n_9349);
  and g19509 (n10418, n10253, n10417);
  not g19510 (n_9350, n10253);
  not g19511 (n_9351, n10417);
  and g19512 (n10419, n_9350, n_9351);
  not g19513 (n_9352, n10248);
  not g19514 (n_9353, n10419);
  and g19515 (n10420, n_9352, n_9353);
  not g19516 (n_9354, n10418);
  and g19517 (n10421, n_9354, n10420);
  not g19518 (n_9355, n10421);
  and g19519 (n10422, n_9352, n_9355);
  and g19520 (n10423, n_9353, n_9355);
  and g19521 (n10424, n_9354, n10423);
  not g19522 (n_9356, n10422);
  not g19523 (n_9357, n10424);
  and g19524 (n10425, n_9356, n_9357);
  not g19525 (n_9358, n10151);
  not g19526 (n_9359, n10425);
  and g19527 (n10426, n_9358, n_9359);
  and g19528 (n10427, n10151, n10425);
  not g19529 (n_9360, n10426);
  not g19530 (n_9361, n10427);
  and g19531 (n10428, n_9360, n_9361);
  not g19532 (n_9362, n10150);
  and g19533 (n10429, n_9362, n10428);
  not g19534 (n_9363, n10428);
  and g19535 (n10430, n10150, n_9363);
  not g19536 (n_9364, n10429);
  not g19537 (n_9365, n10430);
  and g19538 (\asquared[67] , n_9364, n_9365);
  and g19539 (n10432, n_9203, n_9355);
  and g19540 (n10433, n_9133, n_9198);
  and g19541 (n10434, n_9328, n_9348);
  and g19542 (n10435, n10433, n10434);
  not g19543 (n_9366, n10433);
  not g19544 (n_9367, n10434);
  and g19545 (n10436, n_9366, n_9367);
  not g19546 (n_9368, n10435);
  not g19547 (n_9369, n10436);
  and g19548 (n10437, n_9368, n_9369);
  and g19549 (n10438, n_9127, n_9130);
  and g19550 (n10439, \a[48] , \a[53] );
  and g19551 (n10440, \a[14] , n10439);
  and g19552 (n10441, \a[17] , n5888);
  not g19553 (n_9370, n10440);
  not g19554 (n_9371, n10441);
  and g19555 (n10442, n_9370, n_9371);
  and g19556 (n10443, \a[14] , \a[53] );
  and g19557 (n10444, n7325, n10443);
  not g19558 (n_9372, n10444);
  and g19559 (n10445, \a[19] , n_9372);
  not g19560 (n_9373, n10442);
  and g19561 (n10446, n_9373, n10445);
  not g19562 (n_9374, n10446);
  and g19563 (n10447, n_9372, n_9374);
  not g19564 (n_9375, n7325);
  not g19565 (n_9376, n10443);
  and g19566 (n10448, n_9375, n_9376);
  not g19567 (n_9377, n10448);
  and g19568 (n10449, n10447, n_9377);
  and g19569 (n10450, \a[48] , n_9374);
  and g19570 (n10451, \a[19] , n10450);
  not g19571 (n_9378, n10449);
  not g19572 (n_9379, n10451);
  and g19573 (n10452, n_9378, n_9379);
  and g19574 (n10453, n2463, n5344);
  and g19575 (n10454, \a[25] , \a[46] );
  and g19576 (n10455, n9527, n10454);
  not g19577 (n_9380, n10453);
  not g19578 (n_9381, n10455);
  and g19579 (n10456, n_9380, n_9381);
  and g19580 (n10457, \a[21] , \a[46] );
  and g19581 (n10458, \a[26] , \a[41] );
  and g19582 (n10459, n10457, n10458);
  not g19583 (n_9382, n10456);
  not g19584 (n_9383, n10459);
  and g19585 (n10460, n_9382, n_9383);
  not g19586 (n_9384, n10460);
  and g19587 (n10461, \a[42] , n_9384);
  and g19588 (n10462, \a[25] , n10461);
  and g19589 (n10463, n_9383, n_9384);
  not g19590 (n_9385, n10457);
  not g19591 (n_9386, n10458);
  and g19592 (n10464, n_9385, n_9386);
  not g19593 (n_9387, n10464);
  and g19594 (n10465, n10463, n_9387);
  not g19595 (n_9388, n10462);
  not g19596 (n_9389, n10465);
  and g19597 (n10466, n_9388, n_9389);
  not g19598 (n_9390, n10452);
  not g19599 (n_9391, n10466);
  and g19600 (n10467, n_9390, n_9391);
  not g19601 (n_9392, n10467);
  and g19602 (n10468, n_9390, n_9392);
  and g19603 (n10469, n_9391, n_9392);
  not g19604 (n_9393, n10468);
  not g19605 (n_9394, n10469);
  and g19606 (n10470, n_9393, n_9394);
  and g19607 (n10471, \a[27] , \a[40] );
  and g19608 (n10472, \a[28] , \a[39] );
  not g19609 (n_9395, n10471);
  not g19610 (n_9396, n10472);
  and g19611 (n10473, n_9395, n_9396);
  and g19612 (n10474, n2331, n4171);
  not g19613 (n_9397, n10474);
  not g19616 (n_9398, n10473);
  not g19618 (n_9399, n10477);
  and g19619 (n10478, \a[63] , n_9399);
  and g19620 (n10479, \a[4] , n10478);
  and g19621 (n10480, n_9397, n_9399);
  and g19622 (n10481, n_9398, n10480);
  not g19623 (n_9400, n10479);
  not g19624 (n_9401, n10481);
  and g19625 (n10482, n_9400, n_9401);
  not g19626 (n_9402, n10470);
  not g19627 (n_9403, n10482);
  and g19628 (n10483, n_9402, n_9403);
  not g19629 (n_9404, n10483);
  and g19630 (n10484, n_9402, n_9404);
  and g19631 (n10485, n_9403, n_9404);
  not g19632 (n_9405, n10484);
  not g19633 (n_9406, n10485);
  and g19634 (n10486, n_9405, n_9406);
  and g19635 (n10487, \a[5] , \a[62] );
  not g19636 (n_9407, \a[34] );
  not g19637 (n_9408, n10487);
  and g19638 (n10488, n_9407, n_9408);
  and g19639 (n10489, \a[62] , n3664);
  and g19640 (n10490, \a[18] , \a[49] );
  not g19641 (n_9409, n10488);
  not g19642 (n_9410, n10489);
  and g19643 (n10491, n_9409, n_9410);
  and g19644 (n10492, n10490, n10491);
  not g19645 (n_9411, n10492);
  and g19646 (n10493, n_9410, n_9411);
  and g19647 (n10494, n_9409, n10493);
  and g19648 (n10495, n10490, n_9411);
  not g19649 (n_9412, n10494);
  not g19650 (n_9413, n10495);
  and g19651 (n10496, n_9412, n_9413);
  and g19652 (n10497, n3143, n3319);
  and g19653 (n10498, n4136, n4150);
  and g19654 (n10499, n3812, n3828);
  not g19655 (n_9414, n10498);
  not g19656 (n_9415, n10499);
  and g19657 (n10500, n_9414, n_9415);
  not g19658 (n_9416, n10497);
  not g19659 (n_9417, n10500);
  and g19660 (n10501, n_9416, n_9417);
  not g19661 (n_9418, n10501);
  and g19662 (n10502, n4136, n_9418);
  and g19663 (n10503, n_9416, n_9418);
  not g19664 (n_9419, n4150);
  not g19665 (n_9420, n6823);
  and g19666 (n10504, n_9419, n_9420);
  not g19667 (n_9421, n10504);
  and g19668 (n10505, n10503, n_9421);
  not g19669 (n_9422, n10502);
  not g19670 (n_9423, n10505);
  and g19671 (n10506, n_9422, n_9423);
  not g19672 (n_9424, n10496);
  not g19673 (n_9425, n10506);
  and g19674 (n10507, n_9424, n_9425);
  not g19675 (n_9426, n10507);
  and g19676 (n10508, n_9424, n_9426);
  and g19677 (n10509, n_9425, n_9426);
  not g19678 (n_9427, n10508);
  not g19679 (n_9428, n10509);
  and g19680 (n10510, n_9427, n_9428);
  and g19681 (n10511, \a[29] , \a[38] );
  and g19682 (n10512, \a[12] , \a[55] );
  and g19683 (n10513, \a[13] , \a[54] );
  not g19684 (n_9429, n10512);
  not g19685 (n_9430, n10513);
  and g19686 (n10514, n_9429, n_9430);
  and g19687 (n10515, n748, n7701);
  not g19688 (n_9431, n10515);
  and g19689 (n10516, n10511, n_9431);
  not g19690 (n_9432, n10514);
  and g19691 (n10517, n_9432, n10516);
  not g19692 (n_9433, n10517);
  and g19693 (n10518, n10511, n_9433);
  and g19694 (n10519, n_9431, n_9433);
  and g19695 (n10520, n_9432, n10519);
  not g19696 (n_9434, n10518);
  not g19697 (n_9435, n10520);
  and g19698 (n10521, n_9434, n_9435);
  not g19699 (n_9436, n10510);
  not g19700 (n_9437, n10521);
  and g19701 (n10522, n_9436, n_9437);
  not g19702 (n_9438, n10522);
  and g19703 (n10523, n_9436, n_9438);
  and g19704 (n10524, n_9437, n_9438);
  not g19705 (n_9439, n10523);
  not g19706 (n_9440, n10524);
  and g19707 (n10525, n_9439, n_9440);
  and g19708 (n10526, \a[8] , \a[59] );
  and g19709 (n10527, \a[9] , \a[58] );
  not g19710 (n_9441, n10526);
  not g19711 (n_9442, n10527);
  and g19712 (n10528, n_9441, n_9442);
  and g19713 (n10529, n432, n8987);
  and g19714 (n10530, n763, n10089);
  and g19715 (n10531, n380, n9509);
  not g19716 (n_9443, n10530);
  not g19717 (n_9444, n10531);
  and g19718 (n10532, n_9443, n_9444);
  not g19719 (n_9445, n10529);
  not g19720 (n_9446, n10532);
  and g19721 (n10533, n_9445, n_9446);
  not g19722 (n_9447, n10533);
  and g19723 (n10534, n_9445, n_9447);
  not g19724 (n_9448, n10528);
  and g19725 (n10535, n_9448, n10534);
  and g19726 (n10536, \a[60] , n_9447);
  and g19727 (n10537, \a[7] , n10536);
  not g19728 (n_9449, n10535);
  not g19729 (n_9450, n10537);
  and g19730 (n10538, n_9449, n_9450);
  and g19731 (n10539, n1666, n5296);
  and g19732 (n10540, n2115, n4811);
  and g19733 (n10541, n1919, n5713);
  not g19734 (n_9451, n10540);
  not g19735 (n_9452, n10541);
  and g19736 (n10542, n_9451, n_9452);
  not g19737 (n_9453, n10539);
  not g19738 (n_9454, n10542);
  and g19739 (n10543, n_9453, n_9454);
  not g19740 (n_9455, n10543);
  and g19741 (n10544, \a[45] , n_9455);
  and g19742 (n10545, \a[22] , n10544);
  and g19743 (n10546, n_9453, n_9455);
  and g19744 (n10547, \a[23] , \a[44] );
  and g19745 (n10548, \a[24] , \a[43] );
  not g19746 (n_9456, n10547);
  not g19747 (n_9457, n10548);
  and g19748 (n10549, n_9456, n_9457);
  not g19749 (n_9458, n10549);
  and g19750 (n10550, n10546, n_9458);
  not g19751 (n_9459, n10545);
  not g19752 (n_9460, n10550);
  and g19753 (n10551, n_9459, n_9460);
  not g19754 (n_9461, n10538);
  not g19755 (n_9462, n10551);
  and g19756 (n10552, n_9461, n_9462);
  not g19757 (n_9463, n10552);
  and g19758 (n10553, n_9461, n_9463);
  and g19759 (n10554, n_9462, n_9463);
  not g19760 (n_9464, n10553);
  not g19761 (n_9465, n10554);
  and g19762 (n10555, n_9464, n_9465);
  and g19763 (n10556, \a[37] , \a[52] );
  and g19764 (n10557, \a[30] , n10556);
  and g19765 (n10558, \a[15] , n10557);
  and g19766 (n10559, n891, n6968);
  not g19767 (n_9466, n10558);
  not g19768 (n_9467, n10559);
  and g19769 (n10560, n_9466, n_9467);
  and g19770 (n10561, \a[16] , \a[51] );
  and g19771 (n10562, \a[30] , \a[37] );
  and g19772 (n10563, n10561, n10562);
  not g19773 (n_9468, n10560);
  not g19774 (n_9469, n10563);
  and g19775 (n10564, n_9468, n_9469);
  not g19776 (n_9470, n10564);
  and g19777 (n10565, \a[52] , n_9470);
  and g19778 (n10566, \a[15] , n10565);
  not g19779 (n_9471, n10561);
  not g19780 (n_9472, n10562);
  and g19781 (n10567, n_9471, n_9472);
  and g19782 (n10568, n_9469, n_9470);
  not g19783 (n_9473, n10567);
  and g19784 (n10569, n_9473, n10568);
  not g19785 (n_9474, n10566);
  not g19786 (n_9475, n10569);
  and g19787 (n10570, n_9474, n_9475);
  not g19788 (n_9476, n10555);
  not g19789 (n_9477, n10570);
  and g19790 (n10571, n_9476, n_9477);
  not g19791 (n_9478, n10571);
  and g19792 (n10572, n_9476, n_9478);
  and g19793 (n10573, n_9477, n_9478);
  not g19794 (n_9479, n10572);
  not g19795 (n_9480, n10573);
  and g19796 (n10574, n_9479, n_9480);
  not g19797 (n_9481, n10525);
  and g19798 (n10575, n_9481, n10574);
  not g19799 (n_9482, n10574);
  and g19800 (n10576, n10525, n_9482);
  not g19801 (n_9483, n10575);
  not g19802 (n_9484, n10576);
  and g19803 (n10577, n_9483, n_9484);
  not g19804 (n_9485, n10486);
  not g19805 (n_9486, n10577);
  and g19806 (n10578, n_9485, n_9486);
  and g19807 (n10579, n10486, n10577);
  not g19808 (n_9487, n10578);
  not g19809 (n_9488, n10579);
  and g19810 (n10580, n_9487, n_9488);
  not g19811 (n_9489, n10438);
  and g19812 (n10581, n_9489, n10580);
  not g19813 (n_9490, n10580);
  and g19814 (n10582, n10438, n_9490);
  not g19815 (n_9491, n10581);
  not g19816 (n_9492, n10582);
  and g19817 (n10583, n_9491, n_9492);
  and g19818 (n10584, n_9176, n_9180);
  and g19819 (n10585, n_9109, n_9113);
  and g19820 (n10586, n10584, n10585);
  not g19821 (n_9493, n10584);
  not g19822 (n_9494, n10585);
  and g19823 (n10587, n_9493, n_9494);
  not g19824 (n_9495, n10586);
  not g19825 (n_9496, n10587);
  and g19826 (n10588, n_9495, n_9496);
  and g19827 (n10589, n_9168, n_9172);
  not g19828 (n_9497, n10588);
  and g19829 (n10590, n_9497, n10589);
  not g19830 (n_9498, n10589);
  and g19831 (n10591, n10588, n_9498);
  not g19832 (n_9499, n10590);
  not g19833 (n_9500, n10591);
  and g19834 (n10592, n_9499, n_9500);
  and g19835 (n10593, n_9184, n_9187);
  and g19836 (n10594, n_9118, n_9122);
  and g19837 (n10595, n10593, n10594);
  not g19838 (n_9501, n10593);
  not g19839 (n_9502, n10594);
  and g19840 (n10596, n_9501, n_9502);
  not g19841 (n_9503, n10595);
  not g19842 (n_9504, n10596);
  and g19843 (n10597, n_9503, n_9504);
  and g19844 (n10598, n10592, n10597);
  not g19845 (n_9505, n10592);
  not g19846 (n_9506, n10597);
  and g19847 (n10599, n_9505, n_9506);
  not g19848 (n_9507, n10598);
  not g19849 (n_9508, n10599);
  and g19850 (n10600, n_9507, n_9508);
  and g19851 (n10601, n10583, n10600);
  not g19852 (n_9509, n10583);
  not g19853 (n_9510, n10600);
  and g19854 (n10602, n_9509, n_9510);
  not g19855 (n_9511, n10601);
  not g19856 (n_9512, n10602);
  and g19857 (n10603, n_9511, n_9512);
  and g19858 (n10604, n10437, n10603);
  not g19859 (n_9513, n10437);
  not g19860 (n_9514, n10603);
  and g19861 (n10605, n_9513, n_9514);
  and g19862 (n10606, n_9209, n_9354);
  and g19863 (n10607, n_9191, n_9195);
  and g19864 (n10608, n_9338, n_9339);
  not g19865 (n_9515, n10608);
  and g19866 (n10609, n_9344, n_9515);
  and g19867 (n10610, n_9272, n_9284);
  and g19868 (n10611, n_9140, n_9152);
  and g19869 (n10612, n10610, n10611);
  not g19870 (n_9516, n10610);
  not g19871 (n_9517, n10611);
  and g19872 (n10613, n_9516, n_9517);
  not g19873 (n_9518, n10612);
  not g19874 (n_9519, n10613);
  and g19875 (n10614, n_9518, n_9519);
  and g19876 (n10615, n_9232, n_9247);
  not g19877 (n_9520, n10614);
  and g19878 (n10616, n_9520, n10615);
  not g19879 (n_9521, n10615);
  and g19880 (n10617, n10614, n_9521);
  not g19881 (n_9522, n10616);
  not g19882 (n_9523, n10617);
  and g19883 (n10618, n_9522, n_9523);
  and g19884 (n10619, n10196, n10260);
  not g19885 (n_9524, n10196);
  not g19886 (n_9525, n10260);
  and g19887 (n10620, n_9524, n_9525);
  not g19888 (n_9526, n10619);
  not g19889 (n_9527, n10620);
  and g19890 (n10621, n_9526, n_9527);
  not g19891 (n_9528, n10621);
  and g19892 (n10622, n10277, n_9528);
  not g19893 (n_9529, n10277);
  and g19894 (n10623, n_9529, n10621);
  not g19895 (n_9530, n10622);
  not g19896 (n_9531, n10623);
  and g19897 (n10624, n_9530, n_9531);
  and g19898 (n10625, n10309, n10343);
  not g19899 (n_9532, n10309);
  not g19900 (n_9533, n10343);
  and g19901 (n10626, n_9532, n_9533);
  not g19902 (n_9534, n10625);
  not g19903 (n_9535, n10626);
  and g19904 (n10627, n_9534, n_9535);
  not g19905 (n_9536, n10627);
  and g19906 (n10628, n10327, n_9536);
  not g19907 (n_9537, n10327);
  and g19908 (n10629, n_9537, n10627);
  not g19909 (n_9538, n10628);
  not g19910 (n_9539, n10629);
  and g19911 (n10630, n_9538, n_9539);
  and g19912 (n10631, \a[6] , \a[61] );
  not g19913 (n_9540, n10382);
  and g19914 (n10632, n_9540, n10631);
  not g19915 (n_9541, n10631);
  and g19916 (n10633, n10382, n_9541);
  not g19917 (n_9542, n10632);
  not g19918 (n_9543, n10633);
  and g19919 (n10634, n_9542, n_9543);
  not g19920 (n_9544, n10634);
  and g19921 (n10635, n10370, n_9544);
  not g19922 (n_9545, n10370);
  and g19923 (n10636, n_9545, n10634);
  not g19924 (n_9546, n10635);
  not g19925 (n_9547, n10636);
  and g19926 (n10637, n_9546, n_9547);
  and g19927 (n10638, n10630, n10637);
  not g19928 (n_9548, n10630);
  not g19929 (n_9549, n10637);
  and g19930 (n10639, n_9548, n_9549);
  not g19931 (n_9550, n10638);
  not g19932 (n_9551, n10639);
  and g19933 (n10640, n_9550, n_9551);
  and g19934 (n10641, n10624, n10640);
  not g19935 (n_9552, n10624);
  not g19936 (n_9553, n10640);
  and g19937 (n10642, n_9552, n_9553);
  not g19938 (n_9554, n10641);
  not g19939 (n_9555, n10642);
  and g19940 (n10643, n_9554, n_9555);
  and g19941 (n10644, n10618, n10643);
  not g19942 (n_9556, n10618);
  not g19943 (n_9557, n10643);
  and g19944 (n10645, n_9556, n_9557);
  not g19945 (n_9558, n10644);
  not g19946 (n_9559, n10645);
  and g19947 (n10646, n_9558, n_9559);
  not g19948 (n_9560, n10609);
  and g19949 (n10647, n_9560, n10646);
  not g19950 (n_9561, n10646);
  and g19951 (n10648, n10609, n_9561);
  not g19952 (n_9562, n10647);
  not g19953 (n_9563, n10648);
  and g19954 (n10649, n_9562, n_9563);
  not g19955 (n_9564, n10649);
  and g19956 (n10650, n10607, n_9564);
  not g19957 (n_9565, n10607);
  and g19958 (n10651, n_9565, n10649);
  not g19959 (n_9566, n10650);
  not g19960 (n_9567, n10651);
  and g19961 (n10652, n_9566, n_9567);
  and g19962 (n10653, n10293, n10357);
  not g19963 (n_9568, n10293);
  not g19964 (n_9569, n10357);
  and g19965 (n10654, n_9568, n_9569);
  not g19966 (n_9570, n10653);
  not g19967 (n_9571, n10654);
  and g19968 (n10655, n_9570, n_9571);
  and g19969 (n10656, n8060, n9985);
  and g19970 (n10657, n723, n8200);
  and g19971 (n10658, \a[20] , \a[57] );
  and g19972 (n10659, n7730, n10658);
  not g19973 (n_9572, n10657);
  not g19974 (n_9573, n10659);
  and g19975 (n10660, n_9572, n_9573);
  not g19976 (n_9574, n10656);
  not g19977 (n_9575, n10660);
  and g19978 (n10661, n_9574, n_9575);
  not g19979 (n_9576, n10661);
  and g19980 (n10662, \a[57] , n_9576);
  and g19981 (n10663, \a[10] , n10662);
  and g19982 (n10664, n_9574, n_9576);
  and g19983 (n10665, \a[11] , \a[56] );
  and g19984 (n10666, \a[20] , \a[47] );
  not g19985 (n_9577, n10665);
  not g19986 (n_9578, n10666);
  and g19987 (n10667, n_9577, n_9578);
  not g19988 (n_9579, n10667);
  and g19989 (n10668, n10664, n_9579);
  not g19990 (n_9580, n10663);
  not g19991 (n_9581, n10668);
  and g19992 (n10669, n_9580, n_9581);
  not g19993 (n_9582, n10669);
  and g19994 (n10670, n10655, n_9582);
  not g19995 (n_9583, n10670);
  and g19996 (n10671, n10655, n_9583);
  and g19997 (n10672, n_9582, n_9583);
  not g19998 (n_9584, n10671);
  not g19999 (n_9585, n10672);
  and g20000 (n10673, n_9584, n_9585);
  and g20001 (n10674, n_9303, n_9315);
  and g20002 (n10675, n10673, n10674);
  not g20003 (n_9586, n10673);
  not g20004 (n_9587, n10674);
  and g20005 (n10676, n_9586, n_9587);
  not g20006 (n_9588, n10675);
  not g20007 (n_9589, n10676);
  and g20008 (n10677, n_9588, n_9589);
  and g20009 (n10678, n_9333, n_9337);
  not g20010 (n_9590, n10677);
  and g20011 (n10679, n_9590, n10678);
  not g20012 (n_9591, n10678);
  and g20013 (n10680, n10677, n_9591);
  not g20014 (n_9592, n10679);
  not g20015 (n_9593, n10680);
  and g20016 (n10681, n_9592, n_9593);
  and g20017 (n10682, n_9318, n_9319);
  not g20018 (n_9594, n10682);
  and g20019 (n10683, n_9324, n_9594);
  and g20020 (n10684, n_9158, n_9164);
  and g20021 (n10685, n10683, n10684);
  not g20022 (n_9595, n10683);
  not g20023 (n_9596, n10684);
  and g20024 (n10686, n_9595, n_9596);
  not g20025 (n_9597, n10685);
  not g20026 (n_9598, n10686);
  and g20027 (n10687, n_9597, n_9598);
  and g20028 (n10688, n10681, n10687);
  not g20029 (n_9599, n10681);
  not g20030 (n_9600, n10687);
  and g20031 (n10689, n_9599, n_9600);
  not g20032 (n_9601, n10688);
  not g20033 (n_9602, n10689);
  and g20034 (n10690, n_9601, n_9602);
  and g20035 (n10691, n10652, n10690);
  not g20036 (n_9603, n10652);
  not g20037 (n_9604, n10690);
  and g20038 (n10692, n_9603, n_9604);
  not g20039 (n_9605, n10691);
  not g20040 (n_9606, n10692);
  and g20041 (n10693, n_9605, n_9606);
  not g20042 (n_9607, n10606);
  and g20043 (n10694, n_9607, n10693);
  not g20044 (n_9608, n10693);
  and g20045 (n10695, n10606, n_9608);
  not g20046 (n_9609, n10694);
  not g20047 (n_9610, n10695);
  and g20048 (n10696, n_9609, n_9610);
  not g20049 (n_9611, n10605);
  and g20050 (n10697, n_9611, n10696);
  not g20051 (n_9612, n10604);
  and g20052 (n10698, n_9612, n10697);
  not g20053 (n_9613, n10698);
  and g20054 (n10699, n10696, n_9613);
  and g20055 (n10700, n_9611, n_9613);
  and g20056 (n10701, n_9612, n10700);
  not g20057 (n_9614, n10699);
  not g20058 (n_9615, n10701);
  and g20059 (n10702, n_9614, n_9615);
  not g20060 (n_9616, n10432);
  not g20061 (n_9617, n10702);
  and g20062 (n10703, n_9616, n_9617);
  and g20063 (n10704, n10432, n10702);
  not g20064 (n_9618, n10703);
  not g20065 (n_9619, n10704);
  and g20066 (n10705, n_9618, n_9619);
  and g20067 (n10706, n_9362, n_9361);
  not g20068 (n_9620, n10706);
  and g20069 (n10707, n_9360, n_9620);
  not g20070 (n_9621, n10705);
  and g20071 (n10708, n_9621, n10707);
  not g20072 (n_9622, n10707);
  and g20073 (n10709, n10705, n_9622);
  not g20074 (n_9623, n10708);
  not g20075 (n_9624, n10709);
  and g20076 (\asquared[68] , n_9623, n_9624);
  and g20077 (n10711, n_9369, n_9612);
  and g20078 (n10712, n_9558, n_9562);
  and g20079 (n10713, n_9481, n_9482);
  not g20080 (n_9625, n10713);
  and g20081 (n10714, n_9487, n_9625);
  and g20082 (n10715, n_9571, n_9583);
  and g20083 (n10716, n_9535, n_9539);
  and g20084 (n10717, n10715, n10716);
  not g20085 (n_9626, n10715);
  not g20086 (n_9627, n10716);
  and g20087 (n10718, n_9626, n_9627);
  not g20088 (n_9628, n10717);
  not g20089 (n_9629, n10718);
  and g20090 (n10719, n_9628, n_9629);
  and g20091 (n10720, n_9463, n_9478);
  not g20092 (n_9630, n10719);
  and g20093 (n10721, n_9630, n10720);
  not g20094 (n_9631, n10720);
  and g20095 (n10722, n10719, n_9631);
  not g20096 (n_9632, n10721);
  not g20097 (n_9633, n10722);
  and g20098 (n10723, n_9632, n_9633);
  and g20099 (n10724, n380, n9512);
  not g20100 (n_9634, n10724);
  and g20101 (n10725, \a[60] , n_9634);
  and g20102 (n10726, \a[8] , n10725);
  and g20103 (n10727, \a[7] , n_9634);
  and g20104 (n10728, \a[61] , n10727);
  not g20105 (n_9635, n10726);
  not g20106 (n_9636, n10728);
  and g20107 (n10729, n_9635, n_9636);
  not g20108 (n_9637, n10493);
  not g20109 (n_9638, n10729);
  and g20110 (n10730, n_9637, n_9638);
  not g20111 (n_9639, n10730);
  and g20112 (n10731, n_9637, n_9639);
  and g20113 (n10732, n_9638, n_9639);
  not g20114 (n_9640, n10731);
  not g20115 (n_9641, n10732);
  and g20116 (n10733, n_9640, n_9641);
  and g20117 (n10734, n_9542, n_9547);
  and g20118 (n10735, n10733, n10734);
  not g20119 (n_9642, n10733);
  not g20120 (n_9643, n10734);
  and g20121 (n10736, n_9642, n_9643);
  not g20122 (n_9644, n10735);
  not g20123 (n_9645, n10736);
  and g20124 (n10737, n_9644, n_9645);
  and g20125 (n10738, n_9527, n_9531);
  not g20126 (n_9646, n10737);
  and g20127 (n10739, n_9646, n10738);
  not g20128 (n_9647, n10738);
  and g20129 (n10740, n10737, n_9647);
  not g20130 (n_9648, n10739);
  not g20131 (n_9649, n10740);
  and g20132 (n10741, n_9648, n_9649);
  and g20133 (n10742, n10723, n10741);
  not g20134 (n_9650, n10723);
  not g20135 (n_9651, n10741);
  and g20136 (n10743, n_9650, n_9651);
  not g20137 (n_9652, n10742);
  not g20138 (n_9653, n10743);
  and g20139 (n10744, n_9652, n_9653);
  not g20140 (n_9654, n10714);
  and g20141 (n10745, n_9654, n10744);
  not g20142 (n_9655, n10744);
  and g20143 (n10746, n10714, n_9655);
  not g20144 (n_9656, n10745);
  not g20145 (n_9657, n10746);
  and g20146 (n10747, n_9656, n_9657);
  not g20147 (n_9658, n10712);
  and g20148 (n10748, n_9658, n10747);
  not g20149 (n_9659, n10748);
  and g20150 (n10749, n_9658, n_9659);
  and g20151 (n10750, n10747, n_9659);
  not g20152 (n_9660, n10749);
  not g20153 (n_9661, n10750);
  and g20154 (n10751, n_9660, n_9661);
  and g20155 (n10752, n_9504, n_9507);
  and g20156 (n10753, n10447, n10463);
  not g20157 (n_9662, n10447);
  not g20158 (n_9663, n10463);
  and g20159 (n10754, n_9662, n_9663);
  not g20160 (n_9664, n10753);
  not g20161 (n_9665, n10754);
  and g20162 (n10755, n_9664, n_9665);
  not g20163 (n_9666, n10755);
  and g20164 (n10756, n10519, n_9666);
  not g20165 (n_9667, n10519);
  and g20166 (n10757, n_9667, n10755);
  not g20167 (n_9668, n10756);
  not g20168 (n_9669, n10757);
  and g20169 (n10758, n_9668, n_9669);
  and g20170 (n10759, n_9392, n_9404);
  and g20171 (n10760, n_9426, n_9438);
  and g20172 (n10761, n10759, n10760);
  not g20173 (n_9670, n10759);
  not g20174 (n_9671, n10760);
  and g20175 (n10762, n_9670, n_9671);
  not g20176 (n_9672, n10761);
  not g20177 (n_9673, n10762);
  and g20178 (n10763, n_9672, n_9673);
  and g20179 (n10764, n10758, n10763);
  not g20180 (n_9674, n10758);
  not g20181 (n_9675, n10763);
  and g20182 (n10765, n_9674, n_9675);
  not g20183 (n_9676, n10764);
  not g20184 (n_9677, n10765);
  and g20185 (n10766, n_9676, n_9677);
  and g20186 (n10767, n_9496, n_9500);
  and g20187 (n10768, n10546, n10664);
  not g20188 (n_9678, n10546);
  not g20189 (n_9679, n10664);
  and g20190 (n10769, n_9678, n_9679);
  not g20191 (n_9680, n10768);
  not g20192 (n_9681, n10769);
  and g20193 (n10770, n_9680, n_9681);
  not g20194 (n_9682, n10770);
  and g20195 (n10771, n10534, n_9682);
  not g20196 (n_9683, n10534);
  and g20197 (n10772, n_9683, n10770);
  not g20198 (n_9684, n10771);
  not g20199 (n_9685, n10772);
  and g20200 (n10773, n_9684, n_9685);
  and g20201 (n10774, n10480, n10503);
  not g20202 (n_9686, n10480);
  not g20203 (n_9687, n10503);
  and g20204 (n10775, n_9686, n_9687);
  not g20205 (n_9688, n10774);
  not g20206 (n_9689, n10775);
  and g20207 (n10776, n_9688, n_9689);
  not g20208 (n_9690, n10776);
  and g20209 (n10777, n10568, n_9690);
  not g20210 (n_9691, n10568);
  and g20211 (n10778, n_9691, n10776);
  not g20212 (n_9692, n10777);
  not g20213 (n_9693, n10778);
  and g20214 (n10779, n_9692, n_9693);
  and g20215 (n10780, n10773, n10779);
  not g20216 (n_9694, n10773);
  not g20217 (n_9695, n10779);
  and g20218 (n10781, n_9694, n_9695);
  not g20219 (n_9696, n10780);
  not g20220 (n_9697, n10781);
  and g20221 (n10782, n_9696, n_9697);
  not g20222 (n_9698, n10767);
  and g20223 (n10783, n_9698, n10782);
  not g20224 (n_9699, n10782);
  and g20225 (n10784, n10767, n_9699);
  not g20226 (n_9700, n10783);
  not g20227 (n_9701, n10784);
  and g20228 (n10785, n_9700, n_9701);
  and g20229 (n10786, n10766, n10785);
  not g20230 (n_9702, n10766);
  not g20231 (n_9703, n10785);
  and g20232 (n10787, n_9702, n_9703);
  not g20233 (n_9704, n10786);
  not g20234 (n_9705, n10787);
  and g20235 (n10788, n_9704, n_9705);
  not g20236 (n_9706, n10752);
  and g20237 (n10789, n_9706, n10788);
  not g20238 (n_9707, n10788);
  and g20239 (n10790, n10752, n_9707);
  not g20240 (n_9708, n10789);
  not g20241 (n_9709, n10790);
  and g20242 (n10791, n_9708, n_9709);
  not g20243 (n_9710, n10751);
  and g20244 (n10792, n_9710, n10791);
  not g20245 (n_9711, n10792);
  and g20246 (n10793, n10791, n_9711);
  and g20247 (n10794, n_9710, n_9711);
  not g20248 (n_9712, n10793);
  not g20249 (n_9713, n10794);
  and g20250 (n10795, n_9712, n_9713);
  not g20251 (n_9714, n10711);
  not g20252 (n_9715, n10795);
  and g20253 (n10796, n_9714, n_9715);
  not g20254 (n_9716, n10796);
  and g20255 (n10797, n_9714, n_9716);
  and g20256 (n10798, n_9715, n_9716);
  not g20257 (n_9717, n10797);
  not g20258 (n_9718, n10798);
  and g20259 (n10799, n_9717, n_9718);
  and g20260 (n10800, n_9567, n_9605);
  and g20261 (n10801, n_9491, n_9511);
  and g20262 (n10802, n_9598, n_9601);
  and g20263 (n10803, n_9550, n_9554);
  and g20264 (n10804, n_9519, n_9523);
  and g20265 (n10805, n10803, n10804);
  not g20266 (n_9719, n10803);
  not g20267 (n_9720, n10804);
  and g20268 (n10806, n_9719, n_9720);
  not g20269 (n_9721, n10805);
  not g20270 (n_9722, n10806);
  and g20271 (n10807, n_9721, n_9722);
  and g20272 (n10808, n_9589, n_9593);
  not g20273 (n_9723, n10807);
  and g20274 (n10809, n_9723, n10808);
  not g20275 (n_9724, n10808);
  and g20276 (n10810, n10807, n_9724);
  not g20277 (n_9725, n10809);
  not g20278 (n_9726, n10810);
  and g20279 (n10811, n_9725, n_9726);
  and g20280 (n10812, n723, n8436);
  and g20281 (n10813, n1076, n8985);
  and g20282 (n10814, n484, n8987);
  not g20283 (n_9727, n10813);
  not g20284 (n_9728, n10814);
  and g20285 (n10815, n_9727, n_9728);
  not g20286 (n_9729, n10812);
  not g20287 (n_9730, n10815);
  and g20288 (n10816, n_9729, n_9730);
  not g20289 (n_9731, n10816);
  and g20290 (n10817, n_9729, n_9731);
  and g20291 (n10818, \a[10] , \a[58] );
  and g20292 (n10819, \a[11] , \a[57] );
  not g20293 (n_9732, n10818);
  not g20294 (n_9733, n10819);
  and g20295 (n10820, n_9732, n_9733);
  not g20296 (n_9734, n10820);
  and g20297 (n10821, n10817, n_9734);
  and g20298 (n10822, \a[59] , n_9731);
  and g20299 (n10823, \a[9] , n10822);
  not g20300 (n_9735, n10821);
  not g20301 (n_9736, n10823);
  and g20302 (n10824, n_9735, n_9736);
  and g20303 (n10825, n2334, n4171);
  and g20304 (n10826, n2041, n3984);
  and g20305 (n10827, n2331, n5413);
  not g20306 (n_9737, n10826);
  not g20307 (n_9738, n10827);
  and g20308 (n10828, n_9737, n_9738);
  not g20309 (n_9739, n10825);
  not g20310 (n_9740, n10828);
  and g20311 (n10829, n_9739, n_9740);
  not g20312 (n_9741, n10829);
  and g20313 (n10830, \a[41] , n_9741);
  and g20314 (n10831, \a[27] , n10830);
  and g20315 (n10832, \a[28] , \a[40] );
  and g20316 (n10833, \a[29] , \a[39] );
  not g20317 (n_9742, n10832);
  not g20318 (n_9743, n10833);
  and g20319 (n10834, n_9742, n_9743);
  and g20320 (n10835, n_9739, n_9741);
  not g20321 (n_9744, n10834);
  and g20322 (n10836, n_9744, n10835);
  not g20323 (n_9745, n10831);
  not g20324 (n_9746, n10836);
  and g20325 (n10837, n_9745, n_9746);
  not g20326 (n_9747, n10824);
  not g20327 (n_9748, n10837);
  and g20328 (n10838, n_9747, n_9748);
  not g20329 (n_9749, n10838);
  and g20330 (n10839, n_9747, n_9749);
  and g20331 (n10840, n_9748, n_9749);
  not g20332 (n_9750, n10839);
  not g20333 (n_9751, n10840);
  and g20334 (n10841, n_9750, n_9751);
  and g20335 (n10842, \a[5] , \a[63] );
  and g20336 (n10843, \a[6] , \a[62] );
  not g20337 (n_9752, n10842);
  not g20338 (n_9753, n10843);
  and g20339 (n10844, n_9752, n_9753);
  and g20340 (n10845, n332, n9792);
  not g20341 (n_9754, n10845);
  not g20344 (n_9755, n10844);
  not g20346 (n_9756, n10848);
  and g20347 (n10849, \a[47] , n_9756);
  and g20348 (n10850, \a[21] , n10849);
  and g20349 (n10851, n_9754, n_9756);
  and g20350 (n10852, n_9755, n10851);
  not g20351 (n_9757, n10850);
  not g20352 (n_9758, n10852);
  and g20353 (n10853, n_9757, n_9758);
  not g20354 (n_9759, n10841);
  not g20355 (n_9760, n10853);
  and g20356 (n10854, n_9759, n_9760);
  not g20357 (n_9761, n10854);
  and g20358 (n10855, n_9759, n_9761);
  and g20359 (n10856, n_9760, n_9761);
  not g20360 (n_9762, n10855);
  not g20361 (n_9763, n10856);
  and g20362 (n10857, n_9762, n_9763);
  and g20363 (n10858, \a[18] , \a[50] );
  and g20364 (n10859, \a[19] , \a[49] );
  not g20365 (n_9764, n10858);
  not g20366 (n_9765, n10859);
  and g20367 (n10860, n_9764, n_9765);
  and g20368 (n10861, n1149, n6325);
  not g20369 (n_9766, n10861);
  and g20370 (n10862, n2972, n_9766);
  not g20371 (n_9767, n10860);
  and g20372 (n10863, n_9767, n10862);
  not g20373 (n_9768, n10863);
  and g20374 (n10864, n_9766, n_9768);
  and g20375 (n10865, n_9767, n10864);
  and g20376 (n10866, n2972, n_9768);
  not g20377 (n_9769, n10865);
  not g20378 (n_9770, n10866);
  and g20379 (n10867, n_9769, n_9770);
  and g20380 (n10868, n3687, n3812);
  and g20381 (n10869, n2488, n3530);
  and g20382 (n10870, n2865, n4565);
  not g20383 (n_9771, n10869);
  not g20384 (n_9772, n10870);
  and g20385 (n10871, n_9771, n_9772);
  not g20386 (n_9773, n10868);
  not g20387 (n_9774, n10871);
  and g20388 (n10872, n_9773, n_9774);
  not g20389 (n_9775, n10872);
  and g20390 (n10873, \a[38] , n_9775);
  and g20391 (n10874, \a[30] , n10873);
  and g20392 (n10875, n_9773, n_9775);
  and g20393 (n10876, \a[31] , \a[37] );
  and g20394 (n10877, \a[32] , \a[36] );
  not g20395 (n_9776, n10876);
  not g20396 (n_9777, n10877);
  and g20397 (n10878, n_9776, n_9777);
  not g20398 (n_9778, n10878);
  and g20399 (n10879, n10875, n_9778);
  not g20400 (n_9779, n10874);
  not g20401 (n_9780, n10879);
  and g20402 (n10880, n_9779, n_9780);
  not g20403 (n_9781, n10867);
  not g20404 (n_9782, n10880);
  and g20405 (n10881, n_9781, n_9782);
  not g20406 (n_9783, n10881);
  and g20407 (n10882, n_9781, n_9783);
  and g20408 (n10883, n_9782, n_9783);
  not g20409 (n_9784, n10882);
  not g20410 (n_9785, n10883);
  and g20411 (n10884, n_9784, n_9785);
  and g20412 (n10885, \a[12] , \a[56] );
  and g20413 (n10886, n7772, n10885);
  and g20414 (n10887, n748, n9161);
  not g20415 (n_9786, n10886);
  not g20416 (n_9787, n10887);
  and g20417 (n10888, n_9786, n_9787);
  and g20418 (n10889, \a[13] , \a[55] );
  and g20419 (n10890, n7772, n10889);
  not g20420 (n_9788, n10888);
  not g20421 (n_9789, n10890);
  and g20422 (n10891, n_9788, n_9789);
  not g20423 (n_9790, n10891);
  and g20424 (n10892, n10885, n_9790);
  and g20425 (n10893, n_9789, n_9790);
  not g20426 (n_9791, n7772);
  not g20427 (n_9792, n10889);
  and g20428 (n10894, n_9791, n_9792);
  not g20429 (n_9793, n10894);
  and g20430 (n10895, n10893, n_9793);
  not g20431 (n_9794, n10892);
  not g20432 (n_9795, n10895);
  and g20433 (n10896, n_9794, n_9795);
  not g20434 (n_9796, n10884);
  not g20435 (n_9797, n10896);
  and g20436 (n10897, n_9796, n_9797);
  not g20437 (n_9798, n10897);
  and g20438 (n10898, n_9796, n_9798);
  and g20439 (n10899, n_9797, n_9798);
  not g20440 (n_9799, n10898);
  not g20441 (n_9800, n10899);
  and g20442 (n10900, n_9799, n_9800);
  and g20443 (n10901, \a[15] , \a[53] );
  and g20444 (n10902, \a[16] , \a[52] );
  not g20445 (n_9801, n10901);
  not g20446 (n_9802, n10902);
  and g20447 (n10903, n_9801, n_9802);
  and g20448 (n10904, n891, n7433);
  and g20449 (n10905, \a[52] , \a[54] );
  and g20450 (n10906, n893, n10905);
  and g20451 (n10907, n895, n7699);
  not g20452 (n_9803, n10906);
  not g20453 (n_9804, n10907);
  and g20454 (n10908, n_9803, n_9804);
  not g20455 (n_9805, n10904);
  not g20456 (n_9806, n10908);
  and g20457 (n10909, n_9805, n_9806);
  not g20458 (n_9807, n10909);
  and g20459 (n10910, n_9805, n_9807);
  not g20460 (n_9808, n10903);
  and g20461 (n10911, n_9808, n10910);
  and g20462 (n10912, \a[54] , n_9807);
  and g20463 (n10913, \a[14] , n10912);
  not g20464 (n_9809, n10911);
  not g20465 (n_9810, n10913);
  and g20466 (n10914, n_9809, n_9810);
  and g20467 (n10915, n1919, n5560);
  not g20468 (n_9811, n10915);
  and g20470 (n10917, \a[23] , \a[45] );
  and g20471 (n10918, \a[22] , \a[46] );
  not g20472 (n_9812, n10917);
  not g20473 (n_9813, n10918);
  and g20474 (n10919, n_9812, n_9813);
  not g20475 (n_9814, n10919);
  not g20478 (n_9815, n10921);
  and g20479 (n10922, \a[48] , n_9815);
  and g20480 (n10923, \a[20] , n10922);
  and g20481 (n10924, n_9811, n_9815);
  and g20482 (n10925, n_9814, n10924);
  not g20483 (n_9816, n10923);
  not g20484 (n_9817, n10925);
  and g20485 (n10926, n_9816, n_9817);
  not g20486 (n_9818, n10914);
  not g20487 (n_9819, n10926);
  and g20488 (n10927, n_9818, n_9819);
  not g20489 (n_9820, n10927);
  and g20490 (n10928, n_9818, n_9820);
  and g20491 (n10929, n_9819, n_9820);
  not g20492 (n_9821, n10928);
  not g20493 (n_9822, n10929);
  and g20494 (n10930, n_9821, n_9822);
  and g20495 (n10931, n2463, n5018);
  and g20496 (n10932, n2301, n4639);
  and g20497 (n10933, n1904, n5296);
  not g20498 (n_9823, n10932);
  not g20499 (n_9824, n10933);
  and g20500 (n10934, n_9823, n_9824);
  not g20501 (n_9825, n10931);
  not g20502 (n_9826, n10934);
  and g20503 (n10935, n_9825, n_9826);
  not g20504 (n_9827, n10935);
  and g20505 (n10936, \a[44] , n_9827);
  and g20506 (n10937, \a[24] , n10936);
  and g20507 (n10938, n_9825, n_9827);
  and g20508 (n10939, \a[25] , \a[43] );
  and g20509 (n10940, \a[26] , \a[42] );
  not g20510 (n_9828, n10939);
  not g20511 (n_9829, n10940);
  and g20512 (n10941, n_9828, n_9829);
  not g20513 (n_9830, n10941);
  and g20514 (n10942, n10938, n_9830);
  not g20515 (n_9831, n10937);
  not g20516 (n_9832, n10942);
  and g20517 (n10943, n_9831, n_9832);
  not g20518 (n_9833, n10930);
  not g20519 (n_9834, n10943);
  and g20520 (n10944, n_9833, n_9834);
  not g20521 (n_9835, n10944);
  and g20522 (n10945, n_9833, n_9835);
  and g20523 (n10946, n_9834, n_9835);
  not g20524 (n_9836, n10945);
  not g20525 (n_9837, n10946);
  and g20526 (n10947, n_9836, n_9837);
  not g20527 (n_9838, n10900);
  and g20528 (n10948, n_9838, n10947);
  not g20529 (n_9839, n10947);
  and g20530 (n10949, n10900, n_9839);
  not g20531 (n_9840, n10948);
  not g20532 (n_9841, n10949);
  and g20533 (n10950, n_9840, n_9841);
  not g20534 (n_9842, n10857);
  not g20535 (n_9843, n10950);
  and g20536 (n10951, n_9842, n_9843);
  and g20537 (n10952, n10857, n10950);
  not g20538 (n_9844, n10951);
  not g20539 (n_9845, n10952);
  and g20540 (n10953, n_9844, n_9845);
  and g20541 (n10954, n10811, n10953);
  not g20542 (n_9846, n10811);
  not g20543 (n_9847, n10953);
  and g20544 (n10955, n_9846, n_9847);
  not g20545 (n_9848, n10954);
  not g20546 (n_9849, n10955);
  and g20547 (n10956, n_9848, n_9849);
  not g20548 (n_9850, n10802);
  and g20549 (n10957, n_9850, n10956);
  not g20550 (n_9851, n10956);
  and g20551 (n10958, n10802, n_9851);
  not g20552 (n_9852, n10957);
  not g20553 (n_9853, n10958);
  and g20554 (n10959, n_9852, n_9853);
  not g20555 (n_9854, n10801);
  and g20556 (n10960, n_9854, n10959);
  not g20557 (n_9855, n10959);
  and g20558 (n10961, n10801, n_9855);
  not g20559 (n_9856, n10960);
  not g20560 (n_9857, n10961);
  and g20561 (n10962, n_9856, n_9857);
  not g20562 (n_9858, n10800);
  and g20563 (n10963, n_9858, n10962);
  not g20564 (n_9859, n10962);
  and g20565 (n10964, n10800, n_9859);
  not g20566 (n_9860, n10963);
  not g20567 (n_9861, n10964);
  and g20568 (n10965, n_9860, n_9861);
  not g20569 (n_9862, n10799);
  not g20570 (n_9863, n10965);
  and g20571 (n10966, n_9862, n_9863);
  and g20572 (n10967, n10799, n10965);
  not g20573 (n_9864, n10966);
  not g20574 (n_9865, n10967);
  and g20575 (n10968, n_9864, n_9865);
  and g20576 (n10969, n_9609, n_9613);
  and g20577 (n10970, n10968, n10969);
  not g20578 (n_9866, n10968);
  not g20579 (n_9867, n10969);
  and g20580 (n10971, n_9866, n_9867);
  not g20581 (n_9868, n10970);
  not g20582 (n_9869, n10971);
  and g20583 (n10972, n_9868, n_9869);
  and g20584 (n10973, n_9619, n_9622);
  not g20585 (n_9870, n10973);
  and g20586 (n10974, n_9618, n_9870);
  not g20587 (n_9871, n10972);
  and g20588 (n10975, n_9871, n10974);
  not g20589 (n_9872, n10974);
  and g20590 (n10976, n10972, n_9872);
  not g20591 (n_9873, n10975);
  not g20592 (n_9874, n10976);
  and g20593 (\asquared[69] , n_9873, n_9874);
  and g20594 (n10978, n_9659, n_9711);
  and g20595 (n10979, n_9848, n_9852);
  and g20596 (n10980, n10978, n10979);
  not g20597 (n_9875, n10978);
  not g20598 (n_9876, n10979);
  and g20599 (n10981, n_9875, n_9876);
  not g20600 (n_9877, n10980);
  not g20601 (n_9878, n10981);
  and g20602 (n10982, n_9877, n_9878);
  and g20603 (n10983, n_9673, n_9676);
  and g20604 (n10984, n1052, n6968);
  and g20605 (n10985, n3134, n6966);
  and g20606 (n10986, n1149, n6564);
  not g20607 (n_9879, n10985);
  not g20608 (n_9880, n10986);
  and g20609 (n10987, n_9879, n_9880);
  not g20610 (n_9881, n10984);
  not g20611 (n_9882, n10987);
  and g20612 (n10988, n_9881, n_9882);
  not g20613 (n_9883, n10988);
  and g20614 (n10989, n_9881, n_9883);
  and g20615 (n10990, \a[17] , \a[52] );
  and g20616 (n10991, \a[18] , \a[51] );
  not g20617 (n_9884, n10990);
  not g20618 (n_9885, n10991);
  and g20619 (n10992, n_9884, n_9885);
  not g20620 (n_9886, n10992);
  and g20621 (n10993, n10989, n_9886);
  and g20622 (n10994, \a[50] , n_9883);
  and g20623 (n10995, \a[19] , n10994);
  not g20624 (n_9887, n10993);
  not g20625 (n_9888, n10995);
  and g20626 (n10996, n_9887, n_9888);
  and g20627 (n10997, n2617, n4171);
  and g20628 (n10998, n3110, n3984);
  and g20629 (n10999, n2334, n5413);
  not g20630 (n_9889, n10998);
  not g20631 (n_9890, n10999);
  and g20632 (n11000, n_9889, n_9890);
  not g20633 (n_9891, n10997);
  not g20634 (n_9892, n11000);
  and g20635 (n11001, n_9891, n_9892);
  not g20636 (n_9893, n11001);
  and g20637 (n11002, \a[41] , n_9893);
  and g20638 (n11003, \a[28] , n11002);
  and g20639 (n11004, n_9891, n_9893);
  and g20640 (n11005, \a[29] , \a[40] );
  and g20641 (n11006, \a[30] , \a[39] );
  not g20642 (n_9894, n11005);
  not g20643 (n_9895, n11006);
  and g20644 (n11007, n_9894, n_9895);
  not g20645 (n_9896, n11007);
  and g20646 (n11008, n11004, n_9896);
  not g20647 (n_9897, n11003);
  not g20648 (n_9898, n11008);
  and g20649 (n11009, n_9897, n_9898);
  not g20650 (n_9899, n10996);
  not g20651 (n_9900, n11009);
  and g20652 (n11010, n_9899, n_9900);
  not g20653 (n_9901, n11010);
  and g20654 (n11011, n_9899, n_9901);
  and g20655 (n11012, n_9900, n_9901);
  not g20656 (n_9902, n11011);
  not g20657 (n_9903, n11012);
  and g20658 (n11013, n_9902, n_9903);
  and g20659 (n11014, n_9681, n_9685);
  and g20660 (n11015, n11013, n11014);
  not g20661 (n_9904, n11013);
  not g20662 (n_9905, n11014);
  and g20663 (n11016, n_9904, n_9905);
  not g20664 (n_9906, n11015);
  not g20665 (n_9907, n11016);
  and g20666 (n11017, n_9906, n_9907);
  and g20667 (n11018, \a[62] , n4133);
  not g20668 (n_9908, n11018);
  and g20669 (n11019, n3319, n_9908);
  not g20670 (n_9909, n11019);
  and g20671 (n11020, n_9908, n_9909);
  and g20672 (n11021, \a[7] , \a[62] );
  not g20673 (n_9910, \a[35] );
  not g20674 (n_9911, n11021);
  and g20675 (n11022, n_9910, n_9911);
  not g20676 (n_9912, n11022);
  and g20677 (n11023, n11020, n_9912);
  and g20678 (n11024, n3319, n_9909);
  not g20679 (n_9913, n11023);
  not g20680 (n_9914, n11024);
  and g20681 (n11025, n_9913, n_9914);
  and g20682 (n11026, n3143, n3687);
  and g20683 (n11027, n2598, n3530);
  and g20684 (n11028, n3812, n4565);
  not g20685 (n_9915, n11027);
  not g20686 (n_9916, n11028);
  and g20687 (n11029, n_9915, n_9916);
  not g20688 (n_9917, n11026);
  not g20689 (n_9918, n11029);
  and g20690 (n11030, n_9917, n_9918);
  not g20691 (n_9919, n11030);
  and g20692 (n11031, \a[38] , n_9919);
  and g20693 (n11032, \a[31] , n11031);
  and g20694 (n11033, n_9917, n_9919);
  and g20695 (n11034, \a[32] , \a[37] );
  not g20696 (n_9920, n7371);
  not g20697 (n_9921, n11034);
  and g20698 (n11035, n_9920, n_9921);
  not g20699 (n_9922, n11035);
  and g20700 (n11036, n11033, n_9922);
  not g20701 (n_9923, n11032);
  not g20702 (n_9924, n11036);
  and g20703 (n11037, n_9923, n_9924);
  not g20704 (n_9925, n11025);
  not g20705 (n_9926, n11037);
  and g20706 (n11038, n_9925, n_9926);
  not g20707 (n_9927, n11038);
  and g20708 (n11039, n_9925, n_9927);
  and g20709 (n11040, n_9926, n_9927);
  not g20710 (n_9928, n11039);
  not g20711 (n_9929, n11040);
  and g20712 (n11041, n_9928, n_9929);
  and g20713 (n11042, n891, n7699);
  and g20714 (n11043, \a[20] , \a[54] );
  and g20715 (n11044, n9806, n11043);
  not g20716 (n_9930, n11042);
  not g20717 (n_9931, n11044);
  and g20718 (n11045, n_9930, n_9931);
  and g20719 (n11046, n6914, n9431);
  not g20720 (n_9932, n11045);
  not g20721 (n_9933, n11046);
  and g20722 (n11047, n_9932, n_9933);
  not g20723 (n_9934, n11047);
  and g20724 (n11048, \a[54] , n_9934);
  and g20725 (n11049, \a[15] , n11048);
  and g20726 (n11050, n_9933, n_9934);
  not g20727 (n_9935, n6914);
  not g20728 (n_9936, n9431);
  and g20729 (n11051, n_9935, n_9936);
  not g20730 (n_9937, n11051);
  and g20731 (n11052, n11050, n_9937);
  not g20732 (n_9938, n11049);
  not g20733 (n_9939, n11052);
  and g20734 (n11053, n_9938, n_9939);
  not g20735 (n_9940, n11041);
  not g20736 (n_9941, n11053);
  and g20737 (n11054, n_9940, n_9941);
  not g20738 (n_9942, n11054);
  and g20739 (n11055, n_9940, n_9942);
  and g20740 (n11056, n_9941, n_9942);
  not g20741 (n_9943, n11055);
  not g20742 (n_9944, n11056);
  and g20743 (n11057, n_9943, n_9944);
  not g20744 (n_9945, n11057);
  and g20745 (n11058, n11017, n_9945);
  not g20746 (n_9946, n11017);
  and g20747 (n11059, n_9946, n11057);
  not g20748 (n_9947, n10983);
  not g20749 (n_9948, n11059);
  and g20750 (n11060, n_9947, n_9948);
  not g20751 (n_9949, n11058);
  and g20752 (n11061, n_9949, n11060);
  not g20753 (n_9950, n11061);
  and g20754 (n11062, n_9947, n_9950);
  and g20755 (n11063, n_9949, n_9950);
  and g20756 (n11064, n_9948, n11063);
  not g20757 (n_9951, n11062);
  not g20758 (n_9952, n11064);
  and g20759 (n11065, n_9951, n_9952);
  and g20760 (n11066, n_9652, n_9656);
  not g20761 (n_9953, n11065);
  not g20762 (n_9954, n11066);
  and g20763 (n11067, n_9953, n_9954);
  not g20764 (n_9955, n11067);
  and g20765 (n11068, n_9953, n_9955);
  and g20766 (n11069, n_9954, n_9955);
  not g20767 (n_9956, n11068);
  not g20768 (n_9957, n11069);
  and g20769 (n11070, n_9956, n_9957);
  and g20770 (n11071, n484, n9509);
  and g20771 (n11072, n378, n8905);
  and g20772 (n11073, n432, n9512);
  not g20773 (n_9958, n11072);
  not g20774 (n_9959, n11073);
  and g20775 (n11074, n_9958, n_9959);
  not g20776 (n_9960, n11071);
  not g20777 (n_9961, n11074);
  and g20778 (n11075, n_9960, n_9961);
  not g20779 (n_9962, n11075);
  and g20780 (n11076, n_9960, n_9962);
  and g20781 (n11077, \a[9] , \a[60] );
  and g20782 (n11078, \a[10] , \a[59] );
  not g20783 (n_9963, n11077);
  not g20784 (n_9964, n11078);
  and g20785 (n11079, n_9963, n_9964);
  not g20786 (n_9965, n11079);
  and g20787 (n11080, n11076, n_9965);
  and g20788 (n11081, \a[61] , n_9962);
  and g20789 (n11082, \a[8] , n11081);
  not g20790 (n_9966, n11080);
  not g20791 (n_9967, n11082);
  and g20792 (n11083, n_9966, n_9967);
  and g20793 (n11084, n1904, n5713);
  and g20794 (n11085, n1547, n7747);
  and g20795 (n11086, n1666, n5560);
  not g20796 (n_9968, n11085);
  not g20797 (n_9969, n11086);
  and g20798 (n11087, n_9968, n_9969);
  not g20799 (n_9970, n11084);
  not g20800 (n_9971, n11087);
  and g20801 (n11088, n_9970, n_9971);
  not g20802 (n_9972, n11088);
  and g20803 (n11089, \a[46] , n_9972);
  and g20804 (n11090, \a[23] , n11089);
  and g20805 (n11091, \a[24] , \a[45] );
  and g20806 (n11092, \a[25] , \a[44] );
  not g20807 (n_9973, n11091);
  not g20808 (n_9974, n11092);
  and g20809 (n11093, n_9973, n_9974);
  and g20810 (n11094, n_9970, n_9972);
  not g20811 (n_9975, n11093);
  and g20812 (n11095, n_9975, n11094);
  not g20813 (n_9976, n11090);
  not g20814 (n_9977, n11095);
  and g20815 (n11096, n_9976, n_9977);
  not g20816 (n_9978, n11083);
  not g20817 (n_9979, n11096);
  and g20818 (n11097, n_9978, n_9979);
  not g20819 (n_9980, n11097);
  and g20820 (n11098, n_9978, n_9980);
  and g20821 (n11099, n_9979, n_9980);
  not g20822 (n_9981, n11098);
  not g20823 (n_9982, n11099);
  and g20824 (n11100, n_9981, n_9982);
  and g20825 (n11101, \a[26] , \a[43] );
  and g20826 (n11102, \a[27] , \a[42] );
  not g20827 (n_9983, n11101);
  not g20828 (n_9984, n11102);
  and g20829 (n11103, n_9983, n_9984);
  and g20830 (n11104, n2227, n5018);
  not g20831 (n_9985, n11104);
  not g20834 (n_9986, n11103);
  not g20836 (n_9987, n11107);
  and g20837 (n11108, \a[63] , n_9987);
  and g20838 (n11109, \a[6] , n11108);
  and g20839 (n11110, n_9985, n_9987);
  and g20840 (n11111, n_9986, n11110);
  not g20841 (n_9988, n11109);
  not g20842 (n_9989, n11111);
  and g20843 (n11112, n_9988, n_9989);
  not g20844 (n_9990, n11100);
  not g20845 (n_9991, n11112);
  and g20846 (n11113, n_9990, n_9991);
  not g20847 (n_9992, n11113);
  and g20848 (n11114, n_9990, n_9992);
  and g20849 (n11115, n_9991, n_9992);
  not g20850 (n_9993, n11114);
  not g20851 (n_9994, n11115);
  and g20852 (n11116, n_9993, n_9994);
  and g20853 (n11117, n_9629, n_9633);
  and g20854 (n11118, n11116, n11117);
  not g20855 (n_9995, n11116);
  not g20856 (n_9996, n11117);
  and g20857 (n11119, n_9995, n_9996);
  not g20858 (n_9997, n11118);
  not g20859 (n_9998, n11119);
  and g20860 (n11120, n_9997, n_9998);
  and g20861 (n11121, n748, n8200);
  and g20862 (n11122, n818, n7942);
  and g20863 (n11123, n602, n8436);
  not g20864 (n_9999, n11122);
  not g20865 (n_10000, n11123);
  and g20866 (n11124, n_9999, n_10000);
  not g20867 (n_10001, n11121);
  not g20868 (n_10002, n11124);
  and g20869 (n11125, n_10001, n_10002);
  not g20870 (n_10003, n11125);
  and g20871 (n11126, \a[58] , n_10003);
  and g20872 (n11127, \a[11] , n11126);
  and g20873 (n11128, n_10001, n_10003);
  and g20874 (n11129, \a[12] , \a[57] );
  and g20875 (n11130, \a[13] , \a[56] );
  not g20876 (n_10004, n11129);
  not g20877 (n_10005, n11130);
  and g20878 (n11131, n_10004, n_10005);
  not g20879 (n_10006, n11131);
  and g20880 (n11132, n11128, n_10006);
  not g20881 (n_10007, n11127);
  not g20882 (n_10008, n11132);
  and g20883 (n11133, n_10007, n_10008);
  and g20884 (n11134, n_9634, n_9639);
  not g20885 (n_10009, n11133);
  and g20886 (n11135, n_10009, n11134);
  not g20887 (n_10010, n11134);
  and g20888 (n11136, n11133, n_10010);
  not g20889 (n_10011, n11135);
  not g20890 (n_10012, n11136);
  and g20891 (n11137, n_10011, n_10012);
  and g20892 (n11138, \a[21] , \a[48] );
  and g20893 (n11139, \a[22] , \a[47] );
  not g20894 (n_10013, n11138);
  not g20895 (n_10014, n11139);
  and g20896 (n11140, n_10013, n_10014);
  and g20897 (n11141, n1574, n6252);
  not g20898 (n_10015, n11141);
  not g20901 (n_10016, n11140);
  not g20903 (n_10017, n11144);
  and g20904 (n11145, \a[55] , n_10017);
  and g20905 (n11146, \a[14] , n11145);
  and g20906 (n11147, n_10015, n_10017);
  and g20907 (n11148, n_10016, n11147);
  not g20908 (n_10018, n11146);
  not g20909 (n_10019, n11148);
  and g20910 (n11149, n_10018, n_10019);
  not g20911 (n_10020, n11137);
  not g20912 (n_10021, n11149);
  and g20913 (n11150, n_10020, n_10021);
  and g20914 (n11151, n11137, n11149);
  not g20915 (n_10022, n11150);
  not g20916 (n_10023, n11151);
  and g20917 (n11152, n_10022, n_10023);
  and g20918 (n11153, n11120, n11152);
  not g20919 (n_10024, n11120);
  not g20920 (n_10025, n11152);
  and g20921 (n11154, n_10024, n_10025);
  not g20922 (n_10026, n11070);
  not g20923 (n_10027, n11154);
  and g20924 (n11155, n_10026, n_10027);
  not g20925 (n_10028, n11153);
  and g20926 (n11156, n_10028, n11155);
  not g20927 (n_10029, n11156);
  and g20928 (n11157, n_10026, n_10029);
  and g20929 (n11158, n_10027, n_10029);
  and g20930 (n11159, n_10028, n11158);
  not g20931 (n_10030, n11157);
  not g20932 (n_10031, n11159);
  and g20933 (n11160, n_10030, n_10031);
  not g20934 (n_10032, n11160);
  and g20935 (n11161, n10982, n_10032);
  not g20936 (n_10033, n10982);
  and g20937 (n11162, n_10033, n11160);
  and g20938 (n11163, n_9856, n_9860);
  and g20939 (n11164, n_9704, n_9708);
  and g20940 (n11165, n_9838, n_9839);
  not g20941 (n_10034, n11165);
  and g20942 (n11166, n_9844, n_10034);
  and g20943 (n11167, n_9696, n_9700);
  and g20944 (n11168, n10893, n10938);
  not g20945 (n_10035, n10893);
  not g20946 (n_10036, n10938);
  and g20947 (n11169, n_10035, n_10036);
  not g20948 (n_10037, n11168);
  not g20949 (n_10038, n11169);
  and g20950 (n11170, n_10037, n_10038);
  not g20951 (n_10039, n11170);
  and g20952 (n11171, n10835, n_10039);
  not g20953 (n_10040, n10835);
  and g20954 (n11172, n_10040, n11170);
  not g20955 (n_10041, n11171);
  not g20956 (n_10042, n11172);
  and g20957 (n11173, n_10041, n_10042);
  and g20958 (n11174, n_9689, n_9693);
  and g20959 (n11175, n_9665, n_9669);
  and g20960 (n11176, n11174, n11175);
  not g20961 (n_10043, n11174);
  not g20962 (n_10044, n11175);
  and g20963 (n11177, n_10043, n_10044);
  not g20964 (n_10045, n11176);
  not g20965 (n_10046, n11177);
  and g20966 (n11178, n_10045, n_10046);
  and g20967 (n11179, n11173, n11178);
  not g20968 (n_10047, n11173);
  not g20969 (n_10048, n11178);
  and g20970 (n11180, n_10047, n_10048);
  not g20971 (n_10049, n11179);
  not g20972 (n_10050, n11180);
  and g20973 (n11181, n_10049, n_10050);
  not g20974 (n_10051, n11167);
  and g20975 (n11182, n_10051, n11181);
  not g20976 (n_10052, n11181);
  and g20977 (n11183, n11167, n_10052);
  not g20978 (n_10053, n11182);
  not g20979 (n_10054, n11183);
  and g20980 (n11184, n_10053, n_10054);
  not g20981 (n_10055, n11166);
  and g20982 (n11185, n_10055, n11184);
  not g20983 (n_10056, n11184);
  and g20984 (n11186, n11166, n_10056);
  not g20985 (n_10057, n11185);
  not g20986 (n_10058, n11186);
  and g20987 (n11187, n_10057, n_10058);
  not g20988 (n_10059, n11187);
  and g20989 (n11188, n11164, n_10059);
  not g20990 (n_10060, n11164);
  and g20991 (n11189, n_10060, n11187);
  not g20992 (n_10061, n11188);
  not g20993 (n_10062, n11189);
  and g20994 (n11190, n_10061, n_10062);
  and g20995 (n11191, n_9722, n_9726);
  and g20996 (n11192, n_9783, n_9798);
  and g20997 (n11193, n_9820, n_9835);
  and g20998 (n11194, n11192, n11193);
  not g20999 (n_10063, n11192);
  not g21000 (n_10064, n11193);
  and g21001 (n11195, n_10063, n_10064);
  not g21002 (n_10065, n11194);
  not g21003 (n_10066, n11195);
  and g21004 (n11196, n_10065, n_10066);
  and g21005 (n11197, n_9645, n_9649);
  not g21006 (n_10067, n11196);
  and g21007 (n11198, n_10067, n11197);
  not g21008 (n_10068, n11197);
  and g21009 (n11199, n11196, n_10068);
  not g21010 (n_10069, n11198);
  not g21011 (n_10070, n11199);
  and g21012 (n11200, n_10069, n_10070);
  and g21013 (n11201, n10817, n10851);
  not g21014 (n_10071, n10817);
  not g21015 (n_10072, n10851);
  and g21016 (n11202, n_10071, n_10072);
  not g21017 (n_10073, n11201);
  not g21018 (n_10074, n11202);
  and g21019 (n11203, n_10073, n_10074);
  not g21020 (n_10075, n11203);
  and g21021 (n11204, n10924, n_10075);
  not g21022 (n_10076, n10924);
  and g21023 (n11205, n_10076, n11203);
  not g21024 (n_10077, n11204);
  not g21025 (n_10078, n11205);
  and g21026 (n11206, n_10077, n_10078);
  and g21027 (n11207, n10864, n10875);
  not g21028 (n_10079, n10864);
  not g21029 (n_10080, n10875);
  and g21030 (n11208, n_10079, n_10080);
  not g21031 (n_10081, n11207);
  not g21032 (n_10082, n11208);
  and g21033 (n11209, n_10081, n_10082);
  not g21034 (n_10083, n11209);
  and g21035 (n11210, n10910, n_10083);
  not g21036 (n_10084, n10910);
  and g21037 (n11211, n_10084, n11209);
  not g21038 (n_10085, n11210);
  not g21039 (n_10086, n11211);
  and g21040 (n11212, n_10085, n_10086);
  and g21041 (n11213, n_9749, n_9761);
  not g21042 (n_10087, n11212);
  and g21043 (n11214, n_10087, n11213);
  not g21044 (n_10088, n11213);
  and g21045 (n11215, n11212, n_10088);
  not g21046 (n_10089, n11214);
  not g21047 (n_10090, n11215);
  and g21048 (n11216, n_10089, n_10090);
  and g21049 (n11217, n11206, n11216);
  not g21050 (n_10091, n11206);
  not g21051 (n_10092, n11216);
  and g21052 (n11218, n_10091, n_10092);
  not g21053 (n_10093, n11217);
  not g21054 (n_10094, n11218);
  and g21055 (n11219, n_10093, n_10094);
  and g21056 (n11220, n11200, n11219);
  not g21057 (n_10095, n11200);
  not g21058 (n_10096, n11219);
  and g21059 (n11221, n_10095, n_10096);
  not g21060 (n_10097, n11220);
  not g21061 (n_10098, n11221);
  and g21062 (n11222, n_10097, n_10098);
  not g21063 (n_10099, n11222);
  and g21064 (n11223, n11191, n_10099);
  not g21065 (n_10100, n11191);
  and g21066 (n11224, n_10100, n11222);
  not g21067 (n_10101, n11223);
  not g21068 (n_10102, n11224);
  and g21069 (n11225, n_10101, n_10102);
  and g21070 (n11226, n11190, n11225);
  not g21071 (n_10103, n11190);
  not g21072 (n_10104, n11225);
  and g21073 (n11227, n_10103, n_10104);
  not g21074 (n_10105, n11226);
  not g21075 (n_10106, n11227);
  and g21076 (n11228, n_10105, n_10106);
  not g21077 (n_10107, n11163);
  and g21078 (n11229, n_10107, n11228);
  not g21079 (n_10108, n11228);
  and g21080 (n11230, n11163, n_10108);
  not g21081 (n_10109, n11229);
  not g21082 (n_10110, n11230);
  and g21083 (n11231, n_10109, n_10110);
  not g21084 (n_10111, n11162);
  and g21085 (n11232, n_10111, n11231);
  not g21086 (n_10112, n11161);
  and g21087 (n11233, n_10112, n11232);
  not g21088 (n_10113, n11233);
  and g21089 (n11234, n11231, n_10113);
  and g21090 (n11235, n_10111, n_10113);
  and g21091 (n11236, n_10112, n11235);
  not g21092 (n_10114, n11234);
  not g21093 (n_10115, n11236);
  and g21094 (n11237, n_10114, n_10115);
  and g21095 (n11238, n_9862, n10965);
  not g21096 (n_10116, n11238);
  and g21097 (n11239, n_9716, n_10116);
  not g21098 (n_10117, n11237);
  not g21099 (n_10118, n11239);
  and g21100 (n11240, n_10117, n_10118);
  and g21101 (n11241, n11237, n11239);
  not g21102 (n_10119, n11240);
  not g21103 (n_10120, n11241);
  and g21104 (n11242, n_10119, n_10120);
  and g21105 (n11243, n_9868, n_9872);
  not g21106 (n_10121, n11243);
  and g21107 (n11244, n_9869, n_10121);
  not g21108 (n_10122, n11242);
  and g21109 (n11245, n_10122, n11244);
  not g21110 (n_10123, n11244);
  and g21111 (n11246, n11242, n_10123);
  not g21112 (n_10124, n11245);
  not g21113 (n_10125, n11246);
  and g21114 (\asquared[70] , n_10124, n_10125);
  and g21115 (n11248, n_10120, n_10123);
  not g21116 (n_10126, n11248);
  and g21117 (n11249, n_10119, n_10126);
  and g21118 (n11250, n_10109, n_10113);
  and g21119 (n11251, n_10062, n_10105);
  and g21120 (n11252, n11004, n11110);
  not g21121 (n_10127, n11004);
  not g21122 (n_10128, n11110);
  and g21123 (n11253, n_10127, n_10128);
  not g21124 (n_10129, n11252);
  not g21125 (n_10130, n11253);
  and g21126 (n11254, n_10129, n_10130);
  not g21127 (n_10131, n11254);
  and g21128 (n11255, n11094, n_10131);
  not g21129 (n_10132, n11094);
  and g21130 (n11256, n_10132, n11254);
  not g21131 (n_10133, n11255);
  not g21132 (n_10134, n11256);
  and g21133 (n11257, n_10133, n_10134);
  and g21134 (n11258, \a[8] , \a[62] );
  not g21135 (n_10135, n11258);
  and g21136 (n11259, n11020, n_10135);
  not g21137 (n_10136, n11020);
  and g21138 (n11260, n_10136, n11258);
  not g21139 (n_10137, n11033);
  not g21140 (n_10138, n11260);
  and g21141 (n11261, n_10137, n_10138);
  not g21142 (n_10139, n11259);
  and g21143 (n11262, n_10139, n11261);
  not g21144 (n_10140, n11262);
  and g21145 (n11263, n_10137, n_10140);
  and g21146 (n11264, n_10138, n_10140);
  and g21147 (n11265, n_10139, n11264);
  not g21148 (n_10141, n11263);
  not g21149 (n_10142, n11265);
  and g21150 (n11266, n_10141, n_10142);
  not g21151 (n_10143, n11266);
  and g21152 (n11267, n11257, n_10143);
  not g21153 (n_10144, n11267);
  and g21154 (n11268, n11257, n_10144);
  and g21155 (n11269, n_10143, n_10144);
  not g21156 (n_10145, n11268);
  not g21157 (n_10146, n11269);
  and g21158 (n11270, n_10145, n_10146);
  and g21159 (n11271, n_9901, n_9907);
  and g21160 (n11272, n11270, n11271);
  not g21161 (n_10147, n11270);
  not g21162 (n_10148, n11271);
  and g21163 (n11273, n_10147, n_10148);
  not g21164 (n_10149, n11272);
  not g21165 (n_10150, n11273);
  and g21166 (n11274, n_10149, n_10150);
  and g21167 (n11275, n_9980, n_9992);
  and g21168 (n11276, n_10009, n_10010);
  not g21169 (n_10151, n11276);
  and g21170 (n11277, n_10022, n_10151);
  and g21171 (n11278, n11275, n11277);
  not g21172 (n_10152, n11275);
  not g21173 (n_10153, n11277);
  and g21174 (n11279, n_10152, n_10153);
  not g21175 (n_10154, n11278);
  not g21176 (n_10155, n11279);
  and g21177 (n11280, n_10154, n_10155);
  and g21178 (n11281, n_9927, n_9942);
  not g21179 (n_10156, n11280);
  and g21180 (n11282, n_10156, n11281);
  not g21181 (n_10157, n11281);
  and g21182 (n11283, n11280, n_10157);
  not g21183 (n_10158, n11282);
  not g21184 (n_10159, n11283);
  and g21185 (n11284, n_10158, n_10159);
  not g21186 (n_10160, n11063);
  and g21187 (n11285, n_10160, n11284);
  not g21188 (n_10161, n11284);
  and g21189 (n11286, n11063, n_10161);
  not g21190 (n_10162, n11285);
  not g21191 (n_10163, n11286);
  and g21192 (n11287, n_10162, n_10163);
  not g21193 (n_10164, n11274);
  not g21194 (n_10165, n11287);
  and g21195 (n11288, n_10164, n_10165);
  and g21196 (n11289, n11274, n11287);
  not g21197 (n_10166, n11251);
  not g21198 (n_10167, n11289);
  and g21199 (n11290, n_10166, n_10167);
  not g21200 (n_10168, n11288);
  and g21201 (n11291, n_10168, n11290);
  not g21202 (n_10169, n11291);
  and g21203 (n11292, n_10166, n_10169);
  and g21204 (n11293, n_10167, n_10169);
  and g21205 (n11294, n_10168, n11293);
  not g21206 (n_10170, n11292);
  not g21207 (n_10171, n11294);
  and g21208 (n11295, n_10170, n_10171);
  and g21209 (n11296, n_10090, n_10093);
  and g21210 (n11297, \a[7] , \a[63] );
  and g21211 (n11298, \a[23] , \a[47] );
  not g21212 (n_10172, n11297);
  not g21213 (n_10173, n11298);
  and g21214 (n11299, n_10172, n_10173);
  and g21215 (n11300, n11297, n11298);
  not g21216 (n_10174, n11300);
  not g21219 (n_10175, n11299);
  not g21221 (n_10176, n11303);
  and g21222 (n11304, n_10174, n_10176);
  and g21223 (n11305, n_10175, n11304);
  and g21224 (n11306, \a[42] , n_10176);
  and g21225 (n11307, \a[28] , n11306);
  not g21226 (n_10177, n11305);
  not g21227 (n_10178, n11307);
  and g21228 (n11308, n_10177, n_10178);
  and g21229 (n11309, n2865, n4171);
  and g21230 (n11310, n3452, n3984);
  and g21231 (n11311, n2617, n5413);
  not g21232 (n_10179, n11310);
  not g21233 (n_10180, n11311);
  and g21234 (n11312, n_10179, n_10180);
  not g21235 (n_10181, n11309);
  not g21236 (n_10182, n11312);
  and g21237 (n11313, n_10181, n_10182);
  not g21238 (n_10183, n11313);
  and g21239 (n11314, \a[41] , n_10183);
  and g21240 (n11315, \a[29] , n11314);
  and g21241 (n11316, n_10181, n_10183);
  and g21242 (n11317, \a[30] , \a[40] );
  and g21243 (n11318, \a[31] , \a[39] );
  not g21244 (n_10184, n11317);
  not g21245 (n_10185, n11318);
  and g21246 (n11319, n_10184, n_10185);
  not g21247 (n_10186, n11319);
  and g21248 (n11320, n11316, n_10186);
  not g21249 (n_10187, n11315);
  not g21250 (n_10188, n11320);
  and g21251 (n11321, n_10187, n_10188);
  not g21252 (n_10189, n11308);
  not g21253 (n_10190, n11321);
  and g21254 (n11322, n_10189, n_10190);
  not g21255 (n_10191, n11322);
  and g21256 (n11323, n_10189, n_10191);
  and g21257 (n11324, n_10190, n_10191);
  not g21258 (n_10192, n11323);
  not g21259 (n_10193, n11324);
  and g21260 (n11325, n_10192, n_10193);
  and g21261 (n11326, n_10082, n_10086);
  and g21262 (n11327, n11325, n11326);
  not g21263 (n_10194, n11325);
  not g21264 (n_10195, n11326);
  and g21265 (n11328, n_10194, n_10195);
  not g21266 (n_10196, n11327);
  not g21267 (n_10197, n11328);
  and g21268 (n11329, n_10196, n_10197);
  and g21269 (n11330, \a[14] , \a[56] );
  and g21270 (n11331, \a[15] , \a[55] );
  not g21271 (n_10198, n11330);
  not g21272 (n_10199, n11331);
  and g21273 (n11332, n_10198, n_10199);
  and g21274 (n11333, n895, n9161);
  not g21275 (n_10200, n11333);
  not g21278 (n_10201, n11332);
  not g21280 (n_10202, n11336);
  and g21281 (n11337, n_10200, n_10202);
  and g21282 (n11338, n_10201, n11337);
  and g21283 (n11339, \a[48] , n_10202);
  and g21284 (n11340, \a[22] , n11339);
  not g21285 (n_10203, n11338);
  not g21286 (n_10204, n11340);
  and g21287 (n11341, n_10203, n_10204);
  and g21288 (n11342, n2227, n5296);
  and g21289 (n11343, n2633, n4811);
  and g21290 (n11344, n2463, n5713);
  not g21291 (n_10205, n11343);
  not g21292 (n_10206, n11344);
  and g21293 (n11345, n_10205, n_10206);
  not g21294 (n_10207, n11342);
  not g21295 (n_10208, n11345);
  and g21296 (n11346, n_10207, n_10208);
  not g21297 (n_10209, n11346);
  and g21298 (n11347, \a[45] , n_10209);
  and g21299 (n11348, \a[25] , n11347);
  and g21300 (n11349, \a[26] , \a[44] );
  and g21301 (n11350, \a[27] , \a[43] );
  not g21302 (n_10210, n11349);
  not g21303 (n_10211, n11350);
  and g21304 (n11351, n_10210, n_10211);
  and g21305 (n11352, n_10207, n_10209);
  not g21306 (n_10212, n11351);
  and g21307 (n11353, n_10212, n11352);
  not g21308 (n_10213, n11348);
  not g21309 (n_10214, n11353);
  and g21310 (n11354, n_10213, n_10214);
  not g21311 (n_10215, n11341);
  not g21312 (n_10216, n11354);
  and g21313 (n11355, n_10215, n_10216);
  not g21314 (n_10217, n11355);
  and g21315 (n11356, n_10215, n_10217);
  and g21316 (n11357, n_10216, n_10217);
  not g21317 (n_10218, n11356);
  not g21318 (n_10219, n11357);
  and g21319 (n11358, n_10218, n_10219);
  and g21320 (n11359, n1490, n6564);
  and g21321 (n11360, n1492, n9934);
  and g21322 (n11361, n1494, n6325);
  not g21323 (n_10220, n11360);
  not g21324 (n_10221, n11361);
  and g21325 (n11362, n_10220, n_10221);
  not g21326 (n_10222, n11359);
  not g21327 (n_10223, n11362);
  and g21328 (n11363, n_10222, n_10223);
  not g21329 (n_10224, n11363);
  and g21330 (n11364, \a[49] , n_10224);
  and g21331 (n11365, \a[21] , n11364);
  and g21332 (n11366, n_10222, n_10224);
  and g21333 (n11367, \a[19] , \a[51] );
  and g21334 (n11368, \a[20] , \a[50] );
  not g21335 (n_10225, n11367);
  not g21336 (n_10226, n11368);
  and g21337 (n11369, n_10225, n_10226);
  not g21338 (n_10227, n11369);
  and g21339 (n11370, n11366, n_10227);
  not g21340 (n_10228, n11365);
  not g21341 (n_10229, n11370);
  and g21342 (n11371, n_10228, n_10229);
  not g21343 (n_10230, n11358);
  not g21344 (n_10231, n11371);
  and g21345 (n11372, n_10230, n_10231);
  not g21346 (n_10232, n11372);
  and g21347 (n11373, n_10230, n_10232);
  and g21348 (n11374, n_10231, n_10232);
  not g21349 (n_10233, n11373);
  not g21350 (n_10234, n11374);
  and g21351 (n11375, n_10233, n_10234);
  not g21352 (n_10235, n11375);
  and g21353 (n11376, n11329, n_10235);
  not g21354 (n_10236, n11329);
  and g21355 (n11377, n_10236, n11375);
  not g21356 (n_10237, n11296);
  not g21357 (n_10238, n11377);
  and g21358 (n11378, n_10237, n_10238);
  not g21359 (n_10239, n11376);
  and g21360 (n11379, n_10239, n11378);
  not g21361 (n_10240, n11379);
  and g21362 (n11380, n_10237, n_10240);
  and g21363 (n11381, n_10239, n_10240);
  and g21364 (n11382, n_10238, n11381);
  not g21365 (n_10241, n11380);
  not g21366 (n_10242, n11382);
  and g21367 (n11383, n_10241, n_10242);
  and g21368 (n11384, n_10053, n_10057);
  and g21369 (n11385, n723, n9509);
  and g21370 (n11386, n1076, n8905);
  and g21371 (n11387, n484, n9512);
  not g21372 (n_10243, n11386);
  not g21373 (n_10244, n11387);
  and g21374 (n11388, n_10243, n_10244);
  not g21375 (n_10245, n11385);
  not g21376 (n_10246, n11388);
  and g21377 (n11389, n_10245, n_10246);
  not g21378 (n_10247, n11389);
  and g21379 (n11390, n_10245, n_10247);
  and g21380 (n11391, \a[10] , \a[60] );
  and g21381 (n11392, \a[11] , \a[59] );
  not g21382 (n_10248, n11391);
  not g21383 (n_10249, n11392);
  and g21384 (n11393, n_10248, n_10249);
  not g21385 (n_10250, n11393);
  and g21386 (n11394, n11390, n_10250);
  and g21387 (n11395, \a[61] , n_10247);
  and g21388 (n11396, \a[9] , n11395);
  not g21389 (n_10251, n11394);
  not g21390 (n_10252, n11396);
  and g21391 (n11397, n_10251, n_10252);
  and g21392 (n11398, n1048, n7699);
  and g21393 (n11399, n1050, n10905);
  and g21394 (n11400, n1052, n7433);
  not g21395 (n_10253, n11399);
  not g21396 (n_10254, n11400);
  and g21397 (n11401, n_10253, n_10254);
  not g21398 (n_10255, n11398);
  not g21399 (n_10256, n11401);
  and g21400 (n11402, n_10255, n_10256);
  not g21401 (n_10257, n11402);
  and g21402 (n11403, n8237, n_10257);
  and g21403 (n11404, n_10255, n_10257);
  and g21404 (n11405, \a[16] , \a[54] );
  not g21405 (n_10258, n9111);
  not g21406 (n_10259, n11405);
  and g21407 (n11406, n_10258, n_10259);
  not g21408 (n_10260, n11406);
  and g21409 (n11407, n11404, n_10260);
  not g21410 (n_10261, n11403);
  not g21411 (n_10262, n11407);
  and g21412 (n11408, n_10261, n_10262);
  not g21413 (n_10263, n11397);
  not g21414 (n_10264, n11408);
  and g21415 (n11409, n_10263, n_10264);
  not g21416 (n_10265, n11409);
  and g21417 (n11410, n_10263, n_10265);
  and g21418 (n11411, n_10264, n_10265);
  not g21419 (n_10266, n11410);
  not g21420 (n_10267, n11411);
  and g21421 (n11412, n_10266, n_10267);
  and g21422 (n11413, n8167, n10301);
  and g21423 (n11414, n748, n8436);
  and g21424 (n11415, \a[24] , \a[58] );
  and g21425 (n11416, n8073, n11415);
  not g21426 (n_10268, n11414);
  not g21427 (n_10269, n11416);
  and g21428 (n11417, n_10268, n_10269);
  not g21429 (n_10270, n11413);
  not g21430 (n_10271, n11417);
  and g21431 (n11418, n_10270, n_10271);
  not g21432 (n_10272, n11418);
  and g21433 (n11419, \a[58] , n_10272);
  and g21434 (n11420, \a[12] , n11419);
  and g21435 (n11421, n_10270, n_10272);
  and g21436 (n11422, \a[13] , \a[57] );
  not g21437 (n_10273, n5231);
  not g21438 (n_10274, n11422);
  and g21439 (n11423, n_10273, n_10274);
  not g21440 (n_10275, n11423);
  and g21441 (n11424, n11421, n_10275);
  not g21442 (n_10276, n11420);
  not g21443 (n_10277, n11424);
  and g21444 (n11425, n_10276, n_10277);
  not g21445 (n_10278, n11412);
  not g21446 (n_10279, n11425);
  and g21447 (n11426, n_10278, n_10279);
  not g21448 (n_10280, n11426);
  and g21449 (n11427, n_10278, n_10280);
  and g21450 (n11428, n_10279, n_10280);
  not g21451 (n_10281, n11427);
  not g21452 (n_10282, n11428);
  and g21453 (n11429, n_10281, n_10282);
  and g21454 (n11430, n10989, n11050);
  not g21455 (n_10283, n10989);
  not g21456 (n_10284, n11050);
  and g21457 (n11431, n_10283, n_10284);
  not g21458 (n_10285, n11430);
  not g21459 (n_10286, n11431);
  and g21460 (n11432, n_10285, n_10286);
  and g21461 (n11433, n3687, n4150);
  and g21462 (n11434, n3143, n4565);
  and g21463 (n11435, \a[34] , \a[38] );
  and g21464 (n11436, n10877, n11435);
  not g21465 (n_10287, n11434);
  not g21466 (n_10288, n11436);
  and g21467 (n11437, n_10287, n_10288);
  not g21468 (n_10289, n11433);
  not g21469 (n_10290, n11437);
  and g21470 (n11438, n_10289, n_10290);
  not g21471 (n_10291, n11438);
  and g21472 (n11439, \a[38] , n_10291);
  and g21473 (n11440, \a[32] , n11439);
  and g21474 (n11441, n_10289, n_10291);
  and g21475 (n11442, \a[33] , \a[37] );
  not g21476 (n_10292, n4595);
  not g21477 (n_10293, n11442);
  and g21478 (n11443, n_10292, n_10293);
  not g21479 (n_10294, n11443);
  and g21480 (n11444, n11441, n_10294);
  not g21481 (n_10295, n11440);
  not g21482 (n_10296, n11444);
  and g21483 (n11445, n_10295, n_10296);
  not g21484 (n_10297, n11445);
  and g21485 (n11446, n11432, n_10297);
  not g21486 (n_10298, n11446);
  and g21487 (n11447, n11432, n_10298);
  and g21488 (n11448, n_10297, n_10298);
  not g21489 (n_10299, n11447);
  not g21490 (n_10300, n11448);
  and g21491 (n11449, n_10299, n_10300);
  and g21492 (n11450, n_10046, n_10049);
  not g21493 (n_10301, n11449);
  not g21494 (n_10302, n11450);
  and g21495 (n11451, n_10301, n_10302);
  and g21496 (n11452, n11449, n11450);
  not g21497 (n_10303, n11451);
  not g21498 (n_10304, n11452);
  and g21499 (n11453, n_10303, n_10304);
  not g21500 (n_10305, n11429);
  and g21501 (n11454, n_10305, n11453);
  not g21502 (n_10306, n11453);
  and g21503 (n11455, n11429, n_10306);
  not g21504 (n_10307, n11454);
  not g21505 (n_10308, n11455);
  and g21506 (n11456, n_10307, n_10308);
  not g21507 (n_10309, n11384);
  and g21508 (n11457, n_10309, n11456);
  not g21509 (n_10310, n11456);
  and g21510 (n11458, n11384, n_10310);
  not g21511 (n_10311, n11457);
  not g21512 (n_10312, n11458);
  and g21513 (n11459, n_10311, n_10312);
  not g21514 (n_10313, n11383);
  and g21515 (n11460, n_10313, n11459);
  not g21516 (n_10314, n11460);
  and g21517 (n11461, n_10313, n_10314);
  and g21518 (n11462, n11459, n_10314);
  not g21519 (n_10315, n11461);
  not g21520 (n_10316, n11462);
  and g21521 (n11463, n_10315, n_10316);
  not g21522 (n_10317, n11295);
  not g21523 (n_10318, n11463);
  and g21524 (n11464, n_10317, n_10318);
  not g21525 (n_10319, n11464);
  and g21526 (n11465, n_10317, n_10319);
  and g21527 (n11466, n_10318, n_10319);
  not g21528 (n_10320, n11465);
  not g21529 (n_10321, n11466);
  and g21530 (n11467, n_10320, n_10321);
  and g21531 (n11468, n_10097, n_10102);
  and g21532 (n11469, n_9998, n_10028);
  and g21533 (n11470, n_10066, n_10070);
  and g21534 (n11471, n11076, n11128);
  not g21535 (n_10322, n11076);
  not g21536 (n_10323, n11128);
  and g21537 (n11472, n_10322, n_10323);
  not g21538 (n_10324, n11471);
  not g21539 (n_10325, n11472);
  and g21540 (n11473, n_10324, n_10325);
  not g21541 (n_10326, n11473);
  and g21542 (n11474, n11147, n_10326);
  not g21543 (n_10327, n11147);
  and g21544 (n11475, n_10327, n11473);
  not g21545 (n_10328, n11474);
  not g21546 (n_10329, n11475);
  and g21547 (n11476, n_10328, n_10329);
  and g21548 (n11477, n_10074, n_10078);
  and g21549 (n11478, n_10038, n_10042);
  and g21550 (n11479, n11477, n11478);
  not g21551 (n_10330, n11477);
  not g21552 (n_10331, n11478);
  and g21553 (n11480, n_10330, n_10331);
  not g21554 (n_10332, n11479);
  not g21555 (n_10333, n11480);
  and g21556 (n11481, n_10332, n_10333);
  and g21557 (n11482, n11476, n11481);
  not g21558 (n_10334, n11476);
  not g21559 (n_10335, n11481);
  and g21560 (n11483, n_10334, n_10335);
  not g21561 (n_10336, n11482);
  not g21562 (n_10337, n11483);
  and g21563 (n11484, n_10336, n_10337);
  not g21564 (n_10338, n11470);
  and g21565 (n11485, n_10338, n11484);
  not g21566 (n_10339, n11485);
  and g21567 (n11486, n_10338, n_10339);
  and g21568 (n11487, n11484, n_10339);
  not g21569 (n_10340, n11486);
  not g21570 (n_10341, n11487);
  and g21571 (n11488, n_10340, n_10341);
  not g21572 (n_10342, n11469);
  not g21573 (n_10343, n11488);
  and g21574 (n11489, n_10342, n_10343);
  not g21575 (n_10344, n11489);
  and g21576 (n11490, n_10342, n_10344);
  and g21577 (n11491, n_10343, n_10344);
  not g21578 (n_10345, n11490);
  not g21579 (n_10346, n11491);
  and g21580 (n11492, n_10345, n_10346);
  not g21581 (n_10347, n11468);
  not g21582 (n_10348, n11492);
  and g21583 (n11493, n_10347, n_10348);
  not g21584 (n_10349, n11493);
  and g21585 (n11494, n_10347, n_10349);
  and g21586 (n11495, n_10348, n_10349);
  not g21587 (n_10350, n11494);
  not g21588 (n_10351, n11495);
  and g21589 (n11496, n_10350, n_10351);
  and g21590 (n11497, n_9955, n_10029);
  and g21591 (n11498, n11496, n11497);
  not g21592 (n_10352, n11496);
  not g21593 (n_10353, n11497);
  and g21594 (n11499, n_10352, n_10353);
  not g21595 (n_10354, n11498);
  not g21596 (n_10355, n11499);
  and g21597 (n11500, n_10354, n_10355);
  and g21598 (n11501, n_9878, n_10112);
  not g21599 (n_10356, n11501);
  and g21600 (n11502, n11500, n_10356);
  not g21601 (n_10357, n11502);
  and g21602 (n11503, n11500, n_10357);
  and g21603 (n11504, n_10356, n_10357);
  not g21604 (n_10358, n11503);
  not g21605 (n_10359, n11504);
  and g21606 (n11505, n_10358, n_10359);
  not g21607 (n_10360, n11467);
  not g21608 (n_10361, n11505);
  and g21609 (n11506, n_10360, n_10361);
  and g21610 (n11507, n11467, n_10359);
  and g21611 (n11508, n_10358, n11507);
  not g21612 (n_10362, n11506);
  not g21613 (n_10363, n11508);
  and g21614 (n11509, n_10362, n_10363);
  not g21615 (n_10364, n11509);
  and g21616 (n11510, n11250, n_10364);
  not g21617 (n_10365, n11250);
  and g21618 (n11511, n_10365, n11509);
  not g21619 (n_10366, n11510);
  not g21620 (n_10367, n11511);
  and g21621 (n11512, n_10366, n_10367);
  not g21622 (n_10368, n11512);
  and g21623 (n11513, n11249, n_10368);
  not g21624 (n_10369, n11249);
  and g21625 (n11514, n_10369, n_10366);
  and g21626 (n11515, n_10367, n11514);
  not g21627 (n_10370, n11513);
  not g21628 (n_10371, n11515);
  and g21629 (\asquared[71] , n_10370, n_10371);
  not g21630 (n_10372, n11514);
  and g21631 (n11517, n_10367, n_10372);
  and g21632 (n11518, n_10357, n_10362);
  and g21633 (n11519, n_10311, n_10314);
  and g21634 (n11520, n_10286, n_10298);
  and g21635 (n11521, n11264, n11520);
  not g21636 (n_10373, n11264);
  not g21637 (n_10374, n11520);
  and g21638 (n11522, n_10373, n_10374);
  not g21639 (n_10375, n11521);
  not g21640 (n_10376, n11522);
  and g21641 (n11523, n_10375, n_10376);
  and g21642 (n11524, n_10130, n_10134);
  not g21643 (n_10377, n11523);
  and g21644 (n11525, n_10377, n11524);
  not g21645 (n_10378, n11524);
  and g21646 (n11526, n11523, n_10378);
  not g21647 (n_10379, n11525);
  not g21648 (n_10380, n11526);
  and g21649 (n11527, n_10379, n_10380);
  and g21650 (n11528, n_10144, n_10150);
  not g21651 (n_10381, n11527);
  and g21652 (n11529, n_10381, n11528);
  not g21653 (n_10382, n11528);
  and g21654 (n11530, n11527, n_10382);
  not g21655 (n_10383, n11529);
  not g21656 (n_10384, n11530);
  and g21657 (n11531, n_10383, n_10384);
  and g21658 (n11532, n_10303, n_10307);
  not g21659 (n_10385, n11531);
  and g21660 (n11533, n_10385, n11532);
  not g21661 (n_10386, n11532);
  and g21662 (n11534, n11531, n_10386);
  not g21663 (n_10387, n11533);
  not g21664 (n_10388, n11534);
  and g21665 (n11535, n_10387, n_10388);
  and g21666 (n11536, n_10162, n_10167);
  not g21667 (n_10389, n11536);
  and g21668 (n11537, n11535, n_10389);
  not g21669 (n_10390, n11535);
  and g21670 (n11538, n_10390, n11536);
  not g21671 (n_10391, n11537);
  not g21672 (n_10392, n11538);
  and g21673 (n11539, n_10391, n_10392);
  not g21674 (n_10393, n11539);
  and g21675 (n11540, n11519, n_10393);
  not g21676 (n_10394, n11519);
  and g21677 (n11541, n_10394, n11539);
  not g21678 (n_10395, n11540);
  not g21679 (n_10396, n11541);
  and g21680 (n11542, n_10395, n_10396);
  and g21681 (n11543, n_10169, n_10319);
  not g21682 (n_10397, n11542);
  and g21683 (n11544, n_10397, n11543);
  not g21684 (n_10398, n11543);
  and g21685 (n11545, n11542, n_10398);
  not g21686 (n_10399, n11544);
  not g21687 (n_10400, n11545);
  and g21688 (n11546, n_10399, n_10400);
  and g21689 (n11547, n_10349, n_10355);
  and g21690 (n11548, n_10265, n_10280);
  and g21691 (n11549, n_10325, n_10329);
  and g21692 (n11550, n11548, n11549);
  not g21693 (n_10401, n11548);
  not g21694 (n_10402, n11549);
  and g21695 (n11551, n_10401, n_10402);
  not g21696 (n_10403, n11550);
  not g21697 (n_10404, n11551);
  and g21698 (n11552, n_10403, n_10404);
  and g21699 (n11553, n_10217, n_10232);
  not g21700 (n_10405, n11552);
  and g21701 (n11554, n_10405, n11553);
  not g21702 (n_10406, n11553);
  and g21703 (n11555, n11552, n_10406);
  not g21704 (n_10407, n11554);
  not g21705 (n_10408, n11555);
  and g21706 (n11556, n_10407, n_10408);
  not g21707 (n_10409, n11381);
  and g21708 (n11557, n_10409, n11556);
  not g21709 (n_10410, n11556);
  and g21710 (n11558, n11381, n_10410);
  not g21711 (n_10411, n11557);
  not g21712 (n_10412, n11558);
  and g21713 (n11559, n_10411, n_10412);
  and g21714 (n11560, n_10191, n_10197);
  and g21715 (n11561, n11390, n11421);
  not g21716 (n_10413, n11390);
  not g21717 (n_10414, n11421);
  and g21718 (n11562, n_10413, n_10414);
  not g21719 (n_10415, n11561);
  not g21720 (n_10416, n11562);
  and g21721 (n11563, n_10415, n_10416);
  not g21722 (n_10417, n11563);
  and g21723 (n11564, n11352, n_10417);
  not g21724 (n_10418, n11352);
  and g21725 (n11565, n_10418, n11563);
  not g21726 (n_10419, n11564);
  not g21727 (n_10420, n11565);
  and g21728 (n11566, n_10419, n_10420);
  and g21729 (n11567, n11316, n11337);
  not g21730 (n_10421, n11316);
  not g21731 (n_10422, n11337);
  and g21732 (n11568, n_10421, n_10422);
  not g21733 (n_10423, n11567);
  not g21734 (n_10424, n11568);
  and g21735 (n11569, n_10423, n_10424);
  not g21736 (n_10425, n11569);
  and g21737 (n11570, n11304, n_10425);
  not g21738 (n_10426, n11304);
  and g21739 (n11571, n_10426, n11569);
  not g21740 (n_10427, n11570);
  not g21741 (n_10428, n11571);
  and g21742 (n11572, n_10427, n_10428);
  not g21743 (n_10429, n11566);
  not g21744 (n_10430, n11572);
  and g21745 (n11573, n_10429, n_10430);
  and g21746 (n11574, n11566, n11572);
  not g21747 (n_10431, n11573);
  not g21748 (n_10432, n11574);
  and g21749 (n11575, n_10431, n_10432);
  not g21750 (n_10433, n11560);
  and g21751 (n11576, n_10433, n11575);
  not g21752 (n_10434, n11575);
  and g21753 (n11577, n11560, n_10434);
  not g21754 (n_10435, n11576);
  not g21755 (n_10436, n11577);
  and g21756 (n11578, n_10435, n_10436);
  and g21757 (n11579, n11559, n11578);
  not g21758 (n_10437, n11559);
  not g21759 (n_10438, n11578);
  and g21760 (n11580, n_10437, n_10438);
  not g21761 (n_10439, n11579);
  not g21762 (n_10440, n11580);
  and g21763 (n11581, n_10439, n_10440);
  not g21764 (n_10441, n11547);
  and g21765 (n11582, n_10441, n11581);
  not g21766 (n_10442, n11581);
  and g21767 (n11583, n11547, n_10442);
  not g21768 (n_10443, n11582);
  not g21769 (n_10444, n11583);
  and g21770 (n11584, n_10443, n_10444);
  and g21771 (n11585, n_10339, n_10344);
  and g21772 (n11586, \a[9] , \a[62] );
  not g21773 (n_10445, \a[36] );
  not g21774 (n_10446, n11586);
  and g21775 (n11587, n_10445, n_10446);
  and g21776 (n11588, \a[36] , \a[62] );
  and g21777 (n11589, \a[9] , n11588);
  not g21778 (n_10447, n11589);
  not g21781 (n_10448, n11587);
  not g21783 (n_10449, n11592);
  and g21784 (n11593, n_10447, n_10449);
  and g21785 (n11594, n_10448, n11593);
  and g21786 (n11595, \a[49] , n_10449);
  and g21787 (n11596, \a[22] , n11595);
  not g21788 (n_10450, n11594);
  not g21789 (n_10451, n11596);
  and g21790 (n11597, n_10450, n_10451);
  and g21791 (n11598, n1490, n6968);
  and g21792 (n11599, n1492, n6966);
  and g21793 (n11600, n1494, n6564);
  not g21794 (n_10452, n11599);
  not g21795 (n_10453, n11600);
  and g21796 (n11601, n_10452, n_10453);
  not g21797 (n_10454, n11598);
  not g21798 (n_10455, n11601);
  and g21799 (n11602, n_10454, n_10455);
  not g21800 (n_10456, n11602);
  and g21801 (n11603, \a[50] , n_10456);
  and g21802 (n11604, \a[21] , n11603);
  and g21803 (n11605, \a[19] , \a[52] );
  and g21804 (n11606, \a[20] , \a[51] );
  not g21805 (n_10457, n11605);
  not g21806 (n_10458, n11606);
  and g21807 (n11607, n_10457, n_10458);
  and g21808 (n11608, n_10454, n_10456);
  not g21809 (n_10459, n11607);
  and g21810 (n11609, n_10459, n11608);
  not g21811 (n_10460, n11604);
  not g21812 (n_10461, n11609);
  and g21813 (n11610, n_10460, n_10461);
  not g21814 (n_10462, n11597);
  not g21815 (n_10463, n11610);
  and g21816 (n11611, n_10462, n_10463);
  not g21817 (n_10464, n11611);
  and g21818 (n11612, n_10462, n_10464);
  and g21819 (n11613, n_10463, n_10464);
  not g21820 (n_10465, n11612);
  not g21821 (n_10466, n11613);
  and g21822 (n11614, n_10465, n_10466);
  and g21823 (n11615, \a[34] , \a[37] );
  and g21824 (n11616, n3828, n11615);
  and g21825 (n11617, n3828, n4563);
  and g21826 (n11618, n4150, n4565);
  not g21827 (n_10467, n11617);
  not g21828 (n_10468, n11618);
  and g21829 (n11619, n_10467, n_10468);
  not g21830 (n_10469, n11616);
  not g21831 (n_10470, n11619);
  and g21832 (n11620, n_10469, n_10470);
  not g21833 (n_10471, n11620);
  and g21834 (n11621, n4563, n_10471);
  and g21835 (n11622, n_10469, n_10471);
  not g21836 (n_10472, n3828);
  not g21837 (n_10473, n11615);
  and g21838 (n11623, n_10472, n_10473);
  not g21839 (n_10474, n11623);
  and g21840 (n11624, n11622, n_10474);
  not g21841 (n_10475, n11621);
  not g21842 (n_10476, n11624);
  and g21843 (n11625, n_10475, n_10476);
  not g21844 (n_10477, n11614);
  not g21845 (n_10478, n11625);
  and g21846 (n11626, n_10477, n_10478);
  not g21847 (n_10479, n11626);
  and g21848 (n11627, n_10477, n_10479);
  and g21849 (n11628, n_10478, n_10479);
  not g21850 (n_10480, n11627);
  not g21851 (n_10481, n11628);
  and g21852 (n11629, n_10480, n_10481);
  and g21853 (n11630, n11404, n11441);
  not g21854 (n_10482, n11404);
  not g21855 (n_10483, n11441);
  and g21856 (n11631, n_10482, n_10483);
  not g21857 (n_10484, n11630);
  not g21858 (n_10485, n11631);
  and g21859 (n11632, n_10484, n_10485);
  and g21860 (n11633, n378, n9909);
  and g21861 (n11634, \a[60] , \a[63] );
  and g21862 (n11635, n961, n11634);
  and g21863 (n11636, n723, n9512);
  not g21864 (n_10486, n11635);
  not g21865 (n_10487, n11636);
  and g21866 (n11637, n_10486, n_10487);
  not g21867 (n_10488, n11633);
  not g21868 (n_10489, n11637);
  and g21869 (n11638, n_10488, n_10489);
  not g21870 (n_10490, n11638);
  and g21871 (n11639, \a[60] , n_10490);
  and g21872 (n11640, \a[11] , n11639);
  and g21873 (n11641, \a[8] , \a[63] );
  and g21874 (n11642, \a[10] , \a[61] );
  not g21875 (n_10491, n11641);
  not g21876 (n_10492, n11642);
  and g21877 (n11643, n_10491, n_10492);
  and g21878 (n11644, n_10488, n_10490);
  not g21879 (n_10493, n11643);
  and g21880 (n11645, n_10493, n11644);
  not g21881 (n_10494, n11640);
  not g21882 (n_10495, n11645);
  and g21883 (n11646, n_10494, n_10495);
  not g21884 (n_10496, n11646);
  and g21885 (n11647, n11632, n_10496);
  not g21886 (n_10497, n11647);
  and g21887 (n11648, n11632, n_10497);
  and g21888 (n11649, n_10496, n_10497);
  not g21889 (n_10498, n11648);
  not g21890 (n_10499, n11649);
  and g21891 (n11650, n_10498, n_10499);
  and g21892 (n11651, n_10333, n_10336);
  not g21893 (n_10500, n11650);
  not g21894 (n_10501, n11651);
  and g21895 (n11652, n_10500, n_10501);
  and g21896 (n11653, n11650, n11651);
  not g21897 (n_10502, n11652);
  not g21898 (n_10503, n11653);
  and g21899 (n11654, n_10502, n_10503);
  not g21900 (n_10504, n11629);
  and g21901 (n11655, n_10504, n11654);
  not g21902 (n_10505, n11654);
  and g21903 (n11656, n11629, n_10505);
  not g21904 (n_10506, n11655);
  not g21905 (n_10507, n11656);
  and g21906 (n11657, n_10506, n_10507);
  not g21907 (n_10508, n11585);
  and g21908 (n11658, n_10508, n11657);
  not g21909 (n_10509, n11657);
  and g21910 (n11659, n11585, n_10509);
  not g21911 (n_10510, n11658);
  not g21912 (n_10511, n11659);
  and g21913 (n11660, n_10510, n_10511);
  and g21914 (n11661, n_10155, n_10159);
  and g21915 (n11662, n2334, n5018);
  and g21916 (n11663, n2041, n4639);
  and g21917 (n11664, n2331, n5296);
  not g21918 (n_10512, n11663);
  not g21919 (n_10513, n11664);
  and g21920 (n11665, n_10512, n_10513);
  not g21921 (n_10514, n11662);
  not g21922 (n_10515, n11665);
  and g21923 (n11666, n_10514, n_10515);
  not g21924 (n_10516, n11666);
  and g21925 (n11667, n_10514, n_10516);
  and g21926 (n11668, \a[28] , \a[43] );
  and g21927 (n11669, \a[29] , \a[42] );
  not g21928 (n_10517, n11668);
  not g21929 (n_10518, n11669);
  and g21930 (n11670, n_10517, n_10518);
  not g21931 (n_10519, n11670);
  and g21932 (n11671, n11667, n_10519);
  and g21933 (n11672, \a[44] , n_10516);
  and g21934 (n11673, \a[27] , n11672);
  not g21935 (n_10520, n11671);
  not g21936 (n_10521, n11673);
  and g21937 (n11674, n_10520, n_10521);
  and g21938 (n11675, n3812, n4171);
  and g21939 (n11676, n2488, n3984);
  and g21940 (n11677, n2865, n5413);
  not g21941 (n_10522, n11676);
  not g21942 (n_10523, n11677);
  and g21943 (n11678, n_10522, n_10523);
  not g21944 (n_10524, n11675);
  not g21945 (n_10525, n11678);
  and g21946 (n11679, n_10524, n_10525);
  not g21947 (n_10526, n11679);
  and g21948 (n11680, \a[41] , n_10526);
  and g21949 (n11681, \a[30] , n11680);
  and g21950 (n11682, \a[31] , \a[40] );
  and g21951 (n11683, \a[32] , \a[39] );
  not g21952 (n_10527, n11682);
  not g21953 (n_10528, n11683);
  and g21954 (n11684, n_10527, n_10528);
  and g21955 (n11685, n_10524, n_10526);
  not g21956 (n_10529, n11684);
  and g21957 (n11686, n_10529, n11685);
  not g21958 (n_10530, n11681);
  not g21959 (n_10531, n11686);
  and g21960 (n11687, n_10530, n_10531);
  not g21961 (n_10532, n11674);
  not g21962 (n_10533, n11687);
  and g21963 (n11688, n_10532, n_10533);
  not g21964 (n_10534, n11688);
  and g21965 (n11689, n_10532, n_10534);
  and g21966 (n11690, n_10533, n_10534);
  not g21967 (n_10535, n11689);
  not g21968 (n_10536, n11690);
  and g21969 (n11691, n_10535, n_10536);
  and g21970 (n11692, \a[17] , \a[54] );
  not g21971 (n_10537, n8564);
  not g21972 (n_10538, n11692);
  and g21973 (n11693, n_10537, n_10538);
  and g21974 (n11694, n1052, n7699);
  not g21975 (n_10539, n11694);
  not g21978 (n_10540, n11693);
  not g21980 (n_10541, n11697);
  and g21981 (n11698, \a[48] , n_10541);
  and g21982 (n11699, \a[23] , n11698);
  and g21983 (n11700, n_10539, n_10541);
  and g21984 (n11701, n_10540, n11700);
  not g21985 (n_10542, n11699);
  not g21986 (n_10543, n11701);
  and g21987 (n11702, n_10542, n_10543);
  not g21988 (n_10544, n11691);
  not g21989 (n_10545, n11702);
  and g21990 (n11703, n_10544, n_10545);
  not g21991 (n_10546, n11703);
  and g21992 (n11704, n_10544, n_10546);
  and g21993 (n11705, n_10545, n_10546);
  not g21994 (n_10547, n11704);
  not g21995 (n_10548, n11705);
  and g21996 (n11706, n_10547, n_10548);
  and g21997 (n11707, n748, n8987);
  not g21998 (n_10549, n11707);
  and g21999 (n11708, \a[58] , n_10549);
  and g22000 (n11709, \a[13] , n11708);
  and g22001 (n11710, \a[59] , n_10549);
  and g22002 (n11711, \a[12] , n11710);
  not g22003 (n_10550, n11709);
  not g22004 (n_10551, n11711);
  and g22005 (n11712, n_10550, n_10551);
  not g22006 (n_10552, n11366);
  not g22007 (n_10553, n11712);
  and g22008 (n11713, n_10552, n_10553);
  not g22009 (n_10554, n11713);
  and g22010 (n11714, n_10552, n_10554);
  and g22011 (n11715, n_10553, n_10554);
  not g22012 (n_10555, n11714);
  not g22013 (n_10556, n11715);
  and g22014 (n11716, n_10555, n_10556);
  and g22015 (n11717, n891, n9161);
  and g22016 (n11718, \a[55] , \a[57] );
  and g22017 (n11719, n893, n11718);
  and g22018 (n11720, n895, n8200);
  not g22019 (n_10557, n11719);
  not g22020 (n_10558, n11720);
  and g22021 (n11721, n_10557, n_10558);
  not g22022 (n_10559, n11717);
  not g22023 (n_10560, n11721);
  and g22024 (n11722, n_10559, n_10560);
  not g22025 (n_10561, n11722);
  and g22026 (n11723, n_10559, n_10561);
  and g22027 (n11724, \a[15] , \a[56] );
  and g22028 (n11725, \a[16] , \a[55] );
  not g22029 (n_10562, n11724);
  not g22030 (n_10563, n11725);
  and g22031 (n11726, n_10562, n_10563);
  not g22032 (n_10564, n11726);
  and g22033 (n11727, n11723, n_10564);
  and g22034 (n11728, \a[57] , n_10561);
  and g22035 (n11729, \a[14] , n11728);
  not g22036 (n_10565, n11727);
  not g22037 (n_10566, n11729);
  and g22038 (n11730, n_10565, n_10566);
  and g22039 (n11731, n2463, n5560);
  and g22040 (n11732, n2301, n5250);
  and g22041 (n11733, n1904, n5666);
  not g22042 (n_10567, n11732);
  not g22043 (n_10568, n11733);
  and g22044 (n11734, n_10567, n_10568);
  not g22045 (n_10569, n11731);
  not g22046 (n_10570, n11734);
  and g22047 (n11735, n_10569, n_10570);
  not g22048 (n_10571, n11735);
  and g22049 (n11736, \a[47] , n_10571);
  and g22050 (n11737, \a[24] , n11736);
  and g22051 (n11738, n_10569, n_10571);
  and g22052 (n11739, \a[26] , \a[45] );
  not g22053 (n_10572, n10454);
  not g22054 (n_10573, n11739);
  and g22055 (n11740, n_10572, n_10573);
  not g22056 (n_10574, n11740);
  and g22057 (n11741, n11738, n_10574);
  not g22058 (n_10575, n11737);
  not g22059 (n_10576, n11741);
  and g22060 (n11742, n_10575, n_10576);
  not g22061 (n_10577, n11730);
  not g22062 (n_10578, n11742);
  and g22063 (n11743, n_10577, n_10578);
  not g22064 (n_10579, n11743);
  and g22065 (n11744, n_10577, n_10579);
  and g22066 (n11745, n_10578, n_10579);
  not g22067 (n_10580, n11744);
  not g22068 (n_10581, n11745);
  and g22069 (n11746, n_10580, n_10581);
  not g22070 (n_10582, n11716);
  and g22071 (n11747, n_10582, n11746);
  not g22072 (n_10583, n11746);
  and g22073 (n11748, n11716, n_10583);
  not g22074 (n_10584, n11747);
  not g22075 (n_10585, n11748);
  and g22076 (n11749, n_10584, n_10585);
  not g22077 (n_10586, n11706);
  not g22078 (n_10587, n11749);
  and g22079 (n11750, n_10586, n_10587);
  and g22080 (n11751, n11706, n11749);
  not g22081 (n_10588, n11750);
  not g22082 (n_10589, n11751);
  and g22083 (n11752, n_10588, n_10589);
  not g22084 (n_10590, n11661);
  and g22085 (n11753, n_10590, n11752);
  not g22086 (n_10591, n11752);
  and g22087 (n11754, n11661, n_10591);
  not g22088 (n_10592, n11753);
  not g22089 (n_10593, n11754);
  and g22090 (n11755, n_10592, n_10593);
  and g22091 (n11756, n11660, n11755);
  not g22092 (n_10594, n11660);
  not g22093 (n_10595, n11755);
  and g22094 (n11757, n_10594, n_10595);
  not g22095 (n_10596, n11756);
  not g22096 (n_10597, n11757);
  and g22097 (n11758, n_10596, n_10597);
  and g22098 (n11759, n11584, n11758);
  not g22099 (n_10598, n11584);
  not g22100 (n_10599, n11758);
  and g22101 (n11760, n_10598, n_10599);
  not g22102 (n_10600, n11759);
  not g22103 (n_10601, n11760);
  and g22104 (n11761, n_10600, n_10601);
  not g22105 (n_10602, n11546);
  not g22106 (n_10603, n11761);
  and g22107 (n11762, n_10602, n_10603);
  and g22108 (n11763, n11546, n11761);
  not g22109 (n_10604, n11762);
  not g22110 (n_10605, n11763);
  and g22111 (n11764, n_10604, n_10605);
  not g22112 (n_10606, n11764);
  and g22113 (n11765, n11518, n_10606);
  not g22114 (n_10607, n11518);
  and g22115 (n11766, n_10607, n11764);
  not g22116 (n_10608, n11765);
  not g22117 (n_10609, n11766);
  and g22118 (n11767, n_10608, n_10609);
  not g22119 (n_10610, n11517);
  not g22120 (n_10611, n11767);
  and g22121 (n11768, n_10610, n_10611);
  and g22122 (n11769, n11517, n11767);
  or g22123 (\asquared[72] , n11768, n11769);
  and g22124 (n11771, n_10610, n_10608);
  not g22125 (n_10612, n11771);
  and g22126 (n11772, n_10609, n_10612);
  and g22127 (n11773, n_10510, n_10596);
  and g22128 (n11774, n_10432, n_10435);
  and g22129 (n11775, n_10485, n_10497);
  and g22130 (n11776, n2865, n5344);
  and g22131 (n11777, n3452, n4807);
  and g22132 (n11778, n2617, n5018);
  not g22133 (n_10613, n11777);
  not g22134 (n_10614, n11778);
  and g22135 (n11779, n_10613, n_10614);
  not g22136 (n_10615, n11776);
  not g22137 (n_10616, n11779);
  and g22138 (n11780, n_10615, n_10616);
  not g22139 (n_10617, n11780);
  and g22140 (n11781, \a[43] , n_10617);
  and g22141 (n11782, \a[29] , n11781);
  and g22142 (n11783, \a[30] , \a[42] );
  not g22143 (n_10618, n4959);
  not g22144 (n_10619, n11783);
  and g22145 (n11784, n_10618, n_10619);
  and g22146 (n11785, n_10615, n_10617);
  not g22147 (n_10620, n11784);
  and g22148 (n11786, n_10620, n11785);
  not g22149 (n_10621, n11782);
  not g22150 (n_10622, n11786);
  and g22151 (n11787, n_10621, n_10622);
  not g22152 (n_10623, n11775);
  not g22153 (n_10624, n11787);
  and g22154 (n11788, n_10623, n_10624);
  not g22155 (n_10625, n11788);
  and g22156 (n11789, n_10623, n_10625);
  and g22157 (n11790, n_10624, n_10625);
  not g22158 (n_10626, n11789);
  not g22159 (n_10627, n11790);
  and g22160 (n11791, n_10626, n_10627);
  and g22161 (n11792, n_10424, n_10428);
  and g22162 (n11793, n11791, n11792);
  not g22163 (n_10628, n11791);
  not g22164 (n_10629, n11792);
  and g22165 (n11794, n_10628, n_10629);
  not g22166 (n_10630, n11793);
  not g22167 (n_10631, n11794);
  and g22168 (n11795, n_10630, n_10631);
  not g22169 (n_10632, n11774);
  and g22170 (n11796, n_10632, n11795);
  not g22171 (n_10633, n11795);
  and g22172 (n11797, n11774, n_10633);
  not g22173 (n_10634, n11796);
  not g22174 (n_10635, n11797);
  and g22175 (n11798, n_10634, n_10635);
  and g22176 (n11799, n_10502, n_10506);
  not g22177 (n_10636, n11798);
  and g22178 (n11800, n_10636, n11799);
  not g22179 (n_10637, n11799);
  and g22180 (n11801, n11798, n_10637);
  not g22181 (n_10638, n11800);
  not g22182 (n_10639, n11801);
  and g22183 (n11802, n_10638, n_10639);
  and g22184 (n11803, n_10411, n_10439);
  not g22185 (n_10640, n11803);
  and g22186 (n11804, n11802, n_10640);
  not g22187 (n_10641, n11802);
  and g22188 (n11805, n_10641, n11803);
  not g22189 (n_10642, n11804);
  not g22190 (n_10643, n11805);
  and g22191 (n11806, n_10642, n_10643);
  not g22192 (n_10644, n11806);
  and g22193 (n11807, n11773, n_10644);
  not g22194 (n_10645, n11773);
  and g22195 (n11808, n_10645, n11806);
  not g22196 (n_10646, n11807);
  not g22197 (n_10647, n11808);
  and g22198 (n11809, n_10646, n_10647);
  and g22199 (n11810, n_10443, n_10600);
  not g22200 (n_10648, n11809);
  and g22201 (n11811, n_10648, n11810);
  not g22202 (n_10649, n11810);
  and g22203 (n11812, n11809, n_10649);
  not g22204 (n_10650, n11811);
  not g22205 (n_10651, n11812);
  and g22206 (n11813, n_10650, n_10651);
  and g22207 (n11814, n_10391, n_10396);
  and g22208 (n11815, n_10534, n_10546);
  and g22209 (n11816, n_10416, n_10420);
  and g22210 (n11817, n11815, n11816);
  not g22211 (n_10652, n11815);
  not g22212 (n_10653, n11816);
  and g22213 (n11818, n_10652, n_10653);
  not g22214 (n_10654, n11817);
  not g22215 (n_10655, n11818);
  and g22216 (n11819, n_10654, n_10655);
  and g22217 (n11820, n_10464, n_10479);
  not g22218 (n_10656, n11819);
  and g22219 (n11821, n_10656, n11820);
  not g22220 (n_10657, n11820);
  and g22221 (n11822, n11819, n_10657);
  not g22222 (n_10658, n11821);
  not g22223 (n_10659, n11822);
  and g22224 (n11823, n_10658, n_10659);
  and g22225 (n11824, n_10588, n_10592);
  not g22226 (n_10660, n11823);
  and g22227 (n11825, n_10660, n11824);
  not g22228 (n_10661, n11824);
  and g22229 (n11826, n11823, n_10661);
  not g22230 (n_10662, n11825);
  not g22231 (n_10663, n11826);
  and g22232 (n11827, n_10662, n_10663);
  and g22233 (n11828, n_10582, n_10583);
  not g22234 (n_10664, n11828);
  and g22235 (n11829, n_10579, n_10664);
  and g22236 (n11830, n11667, n11700);
  not g22237 (n_10665, n11667);
  not g22238 (n_10666, n11700);
  and g22239 (n11831, n_10665, n_10666);
  not g22240 (n_10667, n11830);
  not g22241 (n_10668, n11831);
  and g22242 (n11832, n_10667, n_10668);
  not g22243 (n_10669, n11832);
  and g22244 (n11833, n11685, n_10669);
  not g22245 (n_10670, n11685);
  and g22246 (n11834, n_10670, n11832);
  not g22247 (n_10671, n11833);
  not g22248 (n_10672, n11834);
  and g22249 (n11835, n_10671, n_10672);
  and g22250 (n11836, n11593, n11622);
  not g22251 (n_10673, n11593);
  not g22252 (n_10674, n11622);
  and g22253 (n11837, n_10673, n_10674);
  not g22254 (n_10675, n11836);
  not g22255 (n_10676, n11837);
  and g22256 (n11838, n_10675, n_10676);
  not g22257 (n_10677, n11838);
  and g22258 (n11839, n11608, n_10677);
  not g22259 (n_10678, n11608);
  and g22260 (n11840, n_10678, n11838);
  not g22261 (n_10679, n11839);
  not g22262 (n_10680, n11840);
  and g22263 (n11841, n_10679, n_10680);
  and g22264 (n11842, n11835, n11841);
  not g22265 (n_10681, n11835);
  not g22266 (n_10682, n11841);
  and g22267 (n11843, n_10681, n_10682);
  not g22268 (n_10683, n11842);
  not g22269 (n_10684, n11843);
  and g22270 (n11844, n_10683, n_10684);
  not g22271 (n_10685, n11829);
  and g22272 (n11845, n_10685, n11844);
  not g22273 (n_10686, n11844);
  and g22274 (n11846, n11829, n_10686);
  not g22275 (n_10687, n11845);
  not g22276 (n_10688, n11846);
  and g22277 (n11847, n_10687, n_10688);
  and g22278 (n11848, n11827, n11847);
  not g22279 (n_10689, n11827);
  not g22280 (n_10690, n11847);
  and g22281 (n11849, n_10689, n_10690);
  not g22282 (n_10691, n11848);
  not g22283 (n_10692, n11849);
  and g22284 (n11850, n_10691, n_10692);
  not g22285 (n_10693, n11850);
  and g22286 (n11851, n11814, n_10693);
  not g22287 (n_10694, n11814);
  and g22288 (n11852, n_10694, n11850);
  not g22289 (n_10695, n11851);
  not g22290 (n_10696, n11852);
  and g22291 (n11853, n_10695, n_10696);
  and g22292 (n11854, n_10404, n_10408);
  and g22293 (n11855, \a[16] , \a[56] );
  and g22294 (n11856, \a[23] , \a[49] );
  not g22295 (n_10697, n11855);
  not g22296 (n_10698, n11856);
  and g22297 (n11857, n_10697, n_10698);
  and g22298 (n11858, n11855, n11856);
  not g22299 (n_10699, n11858);
  not g22302 (n_10700, n11857);
  not g22304 (n_10701, n11861);
  and g22305 (n11862, n_10699, n_10701);
  and g22306 (n11863, n_10700, n11862);
  and g22307 (n11864, \a[40] , n_10701);
  and g22308 (n11865, \a[32] , n11864);
  not g22309 (n_10702, n11863);
  not g22310 (n_10703, n11865);
  and g22311 (n11866, n_10702, n_10703);
  and g22312 (n11867, \a[21] , \a[51] );
  and g22313 (n11868, \a[22] , \a[50] );
  not g22314 (n_10704, n11867);
  not g22315 (n_10705, n11868);
  and g22316 (n11869, n_10704, n_10705);
  and g22317 (n11870, n1574, n6564);
  not g22318 (n_10706, n11870);
  and g22319 (n11871, n5031, n_10706);
  not g22320 (n_10707, n11869);
  and g22321 (n11872, n_10707, n11871);
  not g22322 (n_10708, n11872);
  and g22323 (n11873, n5031, n_10708);
  and g22324 (n11874, n_10706, n_10708);
  and g22325 (n11875, n_10707, n11874);
  not g22326 (n_10709, n11873);
  not g22327 (n_10710, n11875);
  and g22328 (n11876, n_10709, n_10710);
  not g22329 (n_10711, n11866);
  not g22330 (n_10712, n11876);
  and g22331 (n11877, n_10711, n_10712);
  not g22332 (n_10713, n11877);
  and g22333 (n11878, n_10711, n_10713);
  and g22334 (n11879, n_10712, n_10713);
  not g22335 (n_10714, n11878);
  not g22336 (n_10715, n11879);
  and g22337 (n11880, n_10714, n_10715);
  and g22338 (n11881, \a[17] , \a[55] );
  and g22339 (n11882, n1331, n10905);
  and g22340 (n11883, n1052, n7701);
  and g22341 (n11884, \a[20] , \a[52] );
  and g22342 (n11885, n11881, n11884);
  not g22343 (n_10716, n11883);
  not g22344 (n_10717, n11885);
  and g22345 (n11886, n_10716, n_10717);
  not g22346 (n_10718, n11882);
  not g22347 (n_10719, n11886);
  and g22348 (n11887, n_10718, n_10719);
  not g22349 (n_10720, n11887);
  and g22350 (n11888, n11881, n_10720);
  not g22351 (n_10721, n9036);
  not g22352 (n_10722, n11884);
  and g22353 (n11889, n_10721, n_10722);
  and g22354 (n11890, n_10718, n_10720);
  not g22355 (n_10723, n11889);
  and g22356 (n11891, n_10723, n11890);
  not g22357 (n_10724, n11888);
  not g22358 (n_10725, n11891);
  and g22359 (n11892, n_10724, n_10725);
  not g22360 (n_10726, n11880);
  not g22361 (n_10727, n11892);
  and g22362 (n11893, n_10726, n_10727);
  not g22363 (n_10728, n11893);
  and g22364 (n11894, n_10726, n_10728);
  and g22365 (n11895, n_10727, n_10728);
  not g22366 (n_10729, n11894);
  not g22367 (n_10730, n11895);
  and g22368 (n11896, n_10729, n_10730);
  and g22369 (n11897, n723, n9721);
  and g22370 (n11898, n1076, n9909);
  and g22371 (n11899, n484, n9792);
  not g22372 (n_10731, n11898);
  not g22373 (n_10732, n11899);
  and g22374 (n11900, n_10731, n_10732);
  not g22375 (n_10733, n11897);
  not g22376 (n_10734, n11900);
  and g22377 (n11901, n_10733, n_10734);
  not g22378 (n_10735, n11901);
  and g22379 (n11902, n_10733, n_10735);
  and g22380 (n11903, \a[10] , \a[62] );
  and g22381 (n11904, \a[11] , \a[61] );
  not g22382 (n_10736, n11903);
  not g22383 (n_10737, n11904);
  and g22384 (n11905, n_10736, n_10737);
  not g22385 (n_10738, n11905);
  and g22386 (n11906, n11902, n_10738);
  and g22387 (n11907, \a[63] , n_10735);
  and g22388 (n11908, \a[9] , n11907);
  not g22389 (n_10739, n11906);
  not g22390 (n_10740, n11908);
  and g22391 (n11909, n_10739, n_10740);
  and g22392 (n11910, n_10549, n_10554);
  and g22393 (n11911, \a[24] , \a[48] );
  and g22394 (n11912, \a[25] , \a[47] );
  not g22395 (n_10741, n11911);
  not g22396 (n_10742, n11912);
  and g22397 (n11913, n_10741, n_10742);
  and g22398 (n11914, n1904, n6252);
  not g22399 (n_10743, n11914);
  not g22402 (n_10744, n11913);
  not g22404 (n_10745, n11917);
  and g22405 (n11918, \a[60] , n_10745);
  and g22406 (n11919, \a[12] , n11918);
  and g22407 (n11920, n_10743, n_10745);
  and g22408 (n11921, n_10744, n11920);
  not g22409 (n_10746, n11919);
  not g22410 (n_10747, n11921);
  and g22411 (n11922, n_10746, n_10747);
  not g22412 (n_10748, n11910);
  not g22413 (n_10749, n11922);
  and g22414 (n11923, n_10748, n_10749);
  not g22415 (n_10750, n11923);
  and g22416 (n11924, n_10748, n_10750);
  and g22417 (n11925, n_10749, n_10750);
  not g22418 (n_10751, n11924);
  not g22419 (n_10752, n11925);
  and g22420 (n11926, n_10751, n_10752);
  not g22421 (n_10753, n11909);
  not g22422 (n_10754, n11926);
  and g22423 (n11927, n_10753, n_10754);
  and g22424 (n11928, n11909, n_10752);
  and g22425 (n11929, n_10751, n11928);
  not g22426 (n_10755, n11927);
  not g22427 (n_10756, n11929);
  and g22428 (n11930, n_10755, n_10756);
  not g22429 (n_10757, n11896);
  and g22430 (n11931, n_10757, n11930);
  not g22431 (n_10758, n11930);
  and g22432 (n11932, n11896, n_10758);
  not g22433 (n_10759, n11931);
  not g22434 (n_10760, n11932);
  and g22435 (n11933, n_10759, n_10760);
  not g22436 (n_10761, n11854);
  and g22437 (n11934, n_10761, n11933);
  not g22438 (n_10762, n11933);
  and g22439 (n11935, n11854, n_10762);
  not g22440 (n_10763, n11934);
  not g22441 (n_10764, n11935);
  and g22442 (n11936, n_10763, n_10764);
  and g22443 (n11937, n_10384, n_10388);
  and g22444 (n11938, n11723, n11738);
  not g22445 (n_10765, n11723);
  not g22446 (n_10766, n11738);
  and g22447 (n11939, n_10765, n_10766);
  not g22448 (n_10767, n11938);
  not g22449 (n_10768, n11939);
  and g22450 (n11940, n_10767, n_10768);
  not g22451 (n_10769, n11940);
  and g22452 (n11941, n11644, n_10769);
  not g22453 (n_10770, n11644);
  and g22454 (n11942, n_10770, n11940);
  not g22455 (n_10771, n11941);
  not g22456 (n_10772, n11942);
  and g22457 (n11943, n_10771, n_10772);
  and g22458 (n11944, n_10376, n_10380);
  not g22459 (n_10773, n11943);
  and g22460 (n11945, n_10773, n11944);
  not g22461 (n_10774, n11944);
  and g22462 (n11946, n11943, n_10774);
  not g22463 (n_10775, n11945);
  not g22464 (n_10776, n11946);
  and g22465 (n11947, n_10775, n_10776);
  and g22466 (n11948, n895, n8436);
  and g22467 (n11949, n821, n8985);
  and g22468 (n11950, n745, n8987);
  not g22469 (n_10777, n11949);
  not g22470 (n_10778, n11950);
  and g22471 (n11951, n_10777, n_10778);
  not g22472 (n_10779, n11948);
  not g22473 (n_10780, n11951);
  and g22474 (n11952, n_10779, n_10780);
  not g22475 (n_10781, n11952);
  and g22476 (n11953, n_10779, n_10781);
  and g22477 (n11954, \a[14] , \a[58] );
  and g22478 (n11955, \a[15] , \a[57] );
  not g22479 (n_10782, n11954);
  not g22480 (n_10783, n11955);
  and g22481 (n11956, n_10782, n_10783);
  not g22482 (n_10784, n11956);
  and g22483 (n11957, n11953, n_10784);
  and g22484 (n11958, \a[59] , n_10781);
  and g22485 (n11959, \a[13] , n11958);
  not g22486 (n_10785, n11957);
  not g22487 (n_10786, n11959);
  and g22488 (n11960, n_10785, n_10786);
  and g22489 (n11961, n2331, n5713);
  and g22490 (n11962, n2800, n7747);
  and g22491 (n11963, n2227, n5560);
  not g22492 (n_10787, n11962);
  not g22493 (n_10788, n11963);
  and g22494 (n11964, n_10787, n_10788);
  not g22495 (n_10789, n11961);
  not g22496 (n_10790, n11964);
  and g22497 (n11965, n_10789, n_10790);
  not g22498 (n_10791, n11965);
  and g22499 (n11966, \a[46] , n_10791);
  and g22500 (n11967, \a[26] , n11966);
  and g22501 (n11968, n_10789, n_10791);
  and g22502 (n11969, \a[27] , \a[45] );
  and g22503 (n11970, \a[28] , \a[44] );
  not g22504 (n_10792, n11969);
  not g22505 (n_10793, n11970);
  and g22506 (n11971, n_10792, n_10793);
  not g22507 (n_10794, n11971);
  and g22508 (n11972, n11968, n_10794);
  not g22509 (n_10795, n11967);
  not g22510 (n_10796, n11972);
  and g22511 (n11973, n_10795, n_10796);
  not g22512 (n_10797, n11960);
  not g22513 (n_10798, n11973);
  and g22514 (n11974, n_10797, n_10798);
  not g22515 (n_10799, n11974);
  and g22516 (n11975, n_10797, n_10799);
  and g22517 (n11976, n_10798, n_10799);
  not g22518 (n_10800, n11975);
  not g22519 (n_10801, n11976);
  and g22520 (n11977, n_10800, n_10801);
  and g22521 (n11978, \a[19] , \a[53] );
  and g22522 (n11979, \a[33] , \a[39] );
  not g22523 (n_10802, n11435);
  not g22524 (n_10803, n11979);
  and g22525 (n11980, n_10802, n_10803);
  and g22526 (n11981, n4150, n5083);
  not g22527 (n_10804, n11981);
  and g22528 (n11982, n11978, n_10804);
  not g22529 (n_10805, n11980);
  and g22530 (n11983, n_10805, n11982);
  not g22531 (n_10806, n11983);
  and g22532 (n11984, n11978, n_10806);
  and g22533 (n11985, n_10804, n_10806);
  and g22534 (n11986, n_10805, n11985);
  not g22535 (n_10807, n11984);
  not g22536 (n_10808, n11986);
  and g22537 (n11987, n_10807, n_10808);
  not g22538 (n_10809, n11977);
  not g22539 (n_10810, n11987);
  and g22540 (n11988, n_10809, n_10810);
  not g22541 (n_10811, n11988);
  and g22542 (n11989, n_10809, n_10811);
  and g22543 (n11990, n_10810, n_10811);
  not g22544 (n_10812, n11989);
  not g22545 (n_10813, n11990);
  and g22546 (n11991, n_10812, n_10813);
  not g22547 (n_10814, n11947);
  and g22548 (n11992, n_10814, n11991);
  not g22549 (n_10815, n11991);
  and g22550 (n11993, n11947, n_10815);
  not g22551 (n_10816, n11992);
  not g22552 (n_10817, n11993);
  and g22553 (n11994, n_10816, n_10817);
  not g22554 (n_10818, n11937);
  and g22555 (n11995, n_10818, n11994);
  not g22556 (n_10819, n11995);
  and g22557 (n11996, n_10818, n_10819);
  and g22558 (n11997, n11994, n_10819);
  not g22559 (n_10820, n11996);
  not g22560 (n_10821, n11997);
  and g22561 (n11998, n_10820, n_10821);
  not g22562 (n_10822, n11998);
  and g22563 (n11999, n11936, n_10822);
  not g22564 (n_10823, n11999);
  and g22565 (n12000, n11936, n_10823);
  and g22566 (n12001, n_10822, n_10823);
  not g22567 (n_10824, n12000);
  not g22568 (n_10825, n12001);
  and g22569 (n12002, n_10824, n_10825);
  not g22570 (n_10826, n12002);
  and g22571 (n12003, n11853, n_10826);
  not g22572 (n_10827, n12003);
  and g22573 (n12004, n11853, n_10827);
  and g22574 (n12005, n_10826, n_10827);
  not g22575 (n_10828, n12004);
  not g22576 (n_10829, n12005);
  and g22577 (n12006, n_10828, n_10829);
  not g22578 (n_10830, n11813);
  and g22579 (n12007, n_10830, n12006);
  not g22580 (n_10831, n12006);
  and g22581 (n12008, n11813, n_10831);
  not g22582 (n_10832, n12007);
  not g22583 (n_10833, n12008);
  and g22584 (n12009, n_10832, n_10833);
  and g22585 (n12010, n_10400, n_10605);
  not g22586 (n_10834, n12009);
  and g22587 (n12011, n_10834, n12010);
  not g22588 (n_10835, n12010);
  and g22589 (n12012, n12009, n_10835);
  not g22590 (n_10836, n12011);
  not g22591 (n_10837, n12012);
  and g22592 (n12013, n_10836, n_10837);
  not g22593 (n_10838, n12013);
  and g22594 (n12014, n11772, n_10838);
  not g22595 (n_10839, n11772);
  and g22596 (n12015, n_10839, n_10836);
  and g22597 (n12016, n_10837, n12015);
  not g22598 (n_10840, n12014);
  not g22599 (n_10841, n12016);
  and g22600 (\asquared[73] , n_10840, n_10841);
  not g22601 (n_10842, n12015);
  and g22602 (n12018, n_10837, n_10842);
  and g22603 (n12019, n_10651, n_10833);
  and g22604 (n12020, n_10696, n_10827);
  and g22605 (n12021, n_10819, n_10823);
  and g22606 (n12022, n_10663, n_10691);
  and g22607 (n12023, n_10776, n_10817);
  and g22608 (n12024, n_10768, n_10772);
  and g22609 (n12025, n3143, n5413);
  and g22610 (n12026, n2598, n6453);
  and g22611 (n12027, n3812, n5344);
  not g22612 (n_10843, n12026);
  not g22613 (n_10844, n12027);
  and g22614 (n12028, n_10843, n_10844);
  not g22615 (n_10845, n12025);
  not g22616 (n_10846, n12028);
  and g22617 (n12029, n_10845, n_10846);
  not g22618 (n_10847, n12029);
  and g22619 (n12030, \a[42] , n_10847);
  and g22620 (n12031, \a[31] , n12030);
  and g22621 (n12032, n_10845, n_10847);
  and g22622 (n12033, \a[32] , \a[41] );
  and g22623 (n12034, \a[33] , \a[40] );
  not g22624 (n_10848, n12033);
  not g22625 (n_10849, n12034);
  and g22626 (n12035, n_10848, n_10849);
  not g22627 (n_10850, n12035);
  and g22628 (n12036, n12032, n_10850);
  not g22629 (n_10851, n12031);
  not g22630 (n_10852, n12036);
  and g22631 (n12037, n_10851, n_10852);
  not g22632 (n_10853, n12024);
  not g22633 (n_10854, n12037);
  and g22634 (n12038, n_10853, n_10854);
  not g22635 (n_10855, n12038);
  and g22636 (n12039, n_10853, n_10855);
  and g22637 (n12040, n_10854, n_10855);
  not g22638 (n_10856, n12039);
  not g22639 (n_10857, n12040);
  and g22640 (n12041, n_10856, n_10857);
  and g22641 (n12042, n_10668, n_10672);
  and g22642 (n12043, n12041, n12042);
  not g22643 (n_10858, n12041);
  not g22644 (n_10859, n12042);
  and g22645 (n12044, n_10858, n_10859);
  not g22646 (n_10860, n12043);
  not g22647 (n_10861, n12044);
  and g22648 (n12045, n_10860, n_10861);
  and g22649 (n12046, n_10683, n_10687);
  not g22650 (n_10862, n12046);
  and g22651 (n12047, n12045, n_10862);
  not g22652 (n_10863, n12045);
  and g22653 (n12048, n_10863, n12046);
  not g22654 (n_10864, n12047);
  not g22655 (n_10865, n12048);
  and g22656 (n12049, n_10864, n_10865);
  not g22657 (n_10866, n12023);
  and g22658 (n12050, n_10866, n12049);
  not g22659 (n_10867, n12049);
  and g22660 (n12051, n12023, n_10867);
  not g22661 (n_10868, n12050);
  not g22662 (n_10869, n12051);
  and g22663 (n12052, n_10868, n_10869);
  not g22664 (n_10870, n12022);
  and g22665 (n12053, n_10870, n12052);
  not g22666 (n_10871, n12052);
  and g22667 (n12054, n12022, n_10871);
  not g22668 (n_10872, n12053);
  not g22669 (n_10873, n12054);
  and g22670 (n12055, n_10872, n_10873);
  not g22671 (n_10874, n12021);
  and g22672 (n12056, n_10874, n12055);
  not g22673 (n_10875, n12055);
  and g22674 (n12057, n12021, n_10875);
  not g22675 (n_10876, n12056);
  not g22676 (n_10877, n12057);
  and g22677 (n12058, n_10876, n_10877);
  not g22678 (n_10878, n12058);
  and g22679 (n12059, n12020, n_10878);
  not g22680 (n_10879, n12020);
  and g22681 (n12060, n_10879, n12058);
  not g22682 (n_10880, n12059);
  not g22683 (n_10881, n12060);
  and g22684 (n12061, n_10880, n_10881);
  and g22685 (n12062, n_10642, n_10647);
  and g22686 (n12063, n_10750, n_10755);
  and g22687 (n12064, n_10676, n_10680);
  and g22688 (n12065, n12063, n12064);
  not g22689 (n_10882, n12063);
  not g22690 (n_10883, n12064);
  and g22691 (n12066, n_10882, n_10883);
  not g22692 (n_10884, n12065);
  not g22693 (n_10885, n12066);
  and g22694 (n12067, n_10884, n_10885);
  and g22695 (n12068, n_10799, n_10811);
  not g22696 (n_10886, n12067);
  and g22697 (n12069, n_10886, n12068);
  not g22698 (n_10887, n12068);
  and g22699 (n12070, n12067, n_10887);
  not g22700 (n_10888, n12069);
  not g22701 (n_10889, n12070);
  and g22702 (n12071, n_10888, n_10889);
  and g22703 (n12072, n_10759, n_10763);
  not g22704 (n_10890, n12071);
  and g22705 (n12073, n_10890, n12072);
  not g22706 (n_10891, n12072);
  and g22707 (n12074, n12071, n_10891);
  not g22708 (n_10892, n12073);
  not g22709 (n_10893, n12074);
  and g22710 (n12075, n_10892, n_10893);
  and g22711 (n12076, n_10713, n_10728);
  and g22712 (n12077, \a[13] , \a[60] );
  not g22713 (n_10894, n11874);
  and g22714 (n12078, n_10894, n12077);
  not g22715 (n_10895, n12077);
  and g22716 (n12079, n11874, n_10895);
  not g22717 (n_10896, n12078);
  not g22718 (n_10897, n12079);
  and g22719 (n12080, n_10896, n_10897);
  not g22720 (n_10898, n12080);
  and g22721 (n12081, n11985, n_10898);
  not g22722 (n_10899, n11985);
  and g22723 (n12082, n_10899, n12080);
  not g22724 (n_10900, n12081);
  not g22725 (n_10901, n12082);
  and g22726 (n12083, n_10900, n_10901);
  and g22727 (n12084, n11902, n11920);
  not g22728 (n_10902, n11902);
  not g22729 (n_10903, n11920);
  and g22730 (n12085, n_10902, n_10903);
  not g22731 (n_10904, n12084);
  not g22732 (n_10905, n12085);
  and g22733 (n12086, n_10904, n_10905);
  not g22734 (n_10906, n12086);
  and g22735 (n12087, n11890, n_10906);
  not g22736 (n_10907, n11890);
  and g22737 (n12088, n_10907, n12086);
  not g22738 (n_10908, n12087);
  not g22739 (n_10909, n12088);
  and g22740 (n12089, n_10908, n_10909);
  and g22741 (n12090, n12083, n12089);
  not g22742 (n_10910, n12083);
  not g22743 (n_10911, n12089);
  and g22744 (n12091, n_10910, n_10911);
  not g22745 (n_10912, n12090);
  not g22746 (n_10913, n12091);
  and g22747 (n12092, n_10912, n_10913);
  not g22748 (n_10914, n12076);
  and g22749 (n12093, n_10914, n12092);
  not g22750 (n_10915, n12092);
  and g22751 (n12094, n12076, n_10915);
  not g22752 (n_10916, n12093);
  not g22753 (n_10917, n12094);
  and g22754 (n12095, n_10916, n_10917);
  and g22755 (n12096, n12075, n12095);
  not g22756 (n_10918, n12075);
  not g22757 (n_10919, n12095);
  and g22758 (n12097, n_10918, n_10919);
  not g22759 (n_10920, n12096);
  not g22760 (n_10921, n12097);
  and g22761 (n12098, n_10920, n_10921);
  not g22762 (n_10922, n12098);
  and g22763 (n12099, n12062, n_10922);
  not g22764 (n_10923, n12062);
  and g22765 (n12100, n_10923, n12098);
  not g22766 (n_10924, n12099);
  not g22767 (n_10925, n12100);
  and g22768 (n12101, n_10924, n_10925);
  and g22769 (n12102, \a[11] , \a[62] );
  not g22770 (n_10926, \a[37] );
  not g22771 (n_10927, n12102);
  and g22772 (n12103, n_10926, n_10927);
  and g22773 (n12104, \a[62] , n4561);
  not g22774 (n_10928, n12104);
  not g22777 (n_10929, n12103);
  not g22779 (n_10930, n12107);
  and g22780 (n12108, n_10928, n_10930);
  and g22781 (n12109, n_10929, n12108);
  and g22782 (n12110, \a[50] , n_10930);
  and g22783 (n12111, \a[23] , n12110);
  not g22784 (n_10931, n12109);
  not g22785 (n_10932, n12111);
  and g22786 (n12112, n_10931, n_10932);
  and g22787 (n12113, \a[49] , \a[54] );
  and g22788 (n12114, n1664, n12113);
  and g22789 (n12115, n1149, n7701);
  and g22790 (n12116, n4191, n9801);
  not g22791 (n_10933, n12115);
  not g22792 (n_10934, n12116);
  and g22793 (n12117, n_10933, n_10934);
  not g22794 (n_10935, n12114);
  not g22795 (n_10936, n12117);
  and g22796 (n12118, n_10935, n_10936);
  not g22797 (n_10937, n12118);
  and g22798 (n12119, \a[55] , n_10937);
  and g22799 (n12120, \a[18] , n12119);
  and g22800 (n12121, n_10935, n_10937);
  and g22801 (n12122, \a[24] , \a[49] );
  not g22802 (n_10938, n9039);
  not g22803 (n_10939, n12122);
  and g22804 (n12123, n_10938, n_10939);
  not g22805 (n_10940, n12123);
  and g22806 (n12124, n12121, n_10940);
  not g22807 (n_10941, n12120);
  not g22808 (n_10942, n12124);
  and g22809 (n12125, n_10941, n_10942);
  not g22810 (n_10943, n12112);
  not g22811 (n_10944, n12125);
  and g22812 (n12126, n_10943, n_10944);
  not g22813 (n_10945, n12126);
  and g22814 (n12127, n_10943, n_10945);
  and g22815 (n12128, n_10944, n_10945);
  not g22816 (n_10946, n12127);
  not g22817 (n_10947, n12128);
  and g22818 (n12129, n_10946, n_10947);
  and g22819 (n12130, n1494, n7433);
  and g22820 (n12131, n1693, n7232);
  and g22821 (n12132, n1574, n6968);
  not g22822 (n_10948, n12131);
  not g22823 (n_10949, n12132);
  and g22824 (n12133, n_10948, n_10949);
  not g22825 (n_10950, n12130);
  not g22826 (n_10951, n12133);
  and g22827 (n12134, n_10950, n_10951);
  not g22828 (n_10952, n12134);
  and g22829 (n12135, \a[51] , n_10952);
  and g22830 (n12136, \a[22] , n12135);
  and g22831 (n12137, n_10950, n_10952);
  and g22832 (n12138, \a[20] , \a[53] );
  and g22833 (n12139, \a[21] , \a[52] );
  not g22834 (n_10953, n12138);
  not g22835 (n_10954, n12139);
  and g22836 (n12140, n_10953, n_10954);
  not g22837 (n_10955, n12140);
  and g22838 (n12141, n12137, n_10955);
  not g22839 (n_10956, n12136);
  not g22840 (n_10957, n12141);
  and g22841 (n12142, n_10956, n_10957);
  not g22842 (n_10958, n12129);
  not g22843 (n_10959, n12142);
  and g22844 (n12143, n_10958, n_10959);
  not g22845 (n_10960, n12143);
  and g22846 (n12144, n_10958, n_10960);
  and g22847 (n12145, n_10959, n_10960);
  not g22848 (n_10961, n12144);
  not g22849 (n_10962, n12145);
  and g22850 (n12146, n_10961, n_10962);
  and g22851 (n12147, \a[15] , \a[58] );
  and g22852 (n12148, \a[16] , \a[57] );
  not g22853 (n_10963, n12147);
  not g22854 (n_10964, n12148);
  and g22855 (n12149, n_10963, n_10964);
  and g22856 (n12150, n891, n8436);
  and g22857 (n12151, n893, n8985);
  and g22858 (n12152, n895, n8987);
  not g22859 (n_10965, n12151);
  not g22860 (n_10966, n12152);
  and g22861 (n12153, n_10965, n_10966);
  not g22862 (n_10967, n12150);
  not g22863 (n_10968, n12153);
  and g22864 (n12154, n_10967, n_10968);
  not g22865 (n_10969, n12154);
  and g22866 (n12155, n_10967, n_10969);
  not g22867 (n_10970, n12149);
  and g22868 (n12156, n_10970, n12155);
  and g22869 (n12157, \a[59] , n_10969);
  and g22870 (n12158, \a[14] , n12157);
  not g22871 (n_10971, n12156);
  not g22872 (n_10972, n12158);
  and g22873 (n12159, n_10971, n_10972);
  and g22874 (n12160, \a[26] , \a[47] );
  and g22875 (n12161, \a[27] , \a[46] );
  not g22876 (n_10973, n12160);
  not g22877 (n_10974, n12161);
  and g22878 (n12162, n_10973, n_10974);
  and g22879 (n12163, n2227, n5666);
  not g22880 (n_10975, n12163);
  not g22883 (n_10976, n12162);
  not g22885 (n_10977, n12166);
  and g22886 (n12167, \a[56] , n_10977);
  and g22887 (n12168, \a[17] , n12167);
  and g22888 (n12169, n_10975, n_10977);
  and g22889 (n12170, n_10976, n12169);
  not g22890 (n_10978, n12168);
  not g22891 (n_10979, n12170);
  and g22892 (n12171, n_10978, n_10979);
  not g22893 (n_10980, n11862);
  not g22894 (n_10981, n12171);
  and g22895 (n12172, n_10980, n_10981);
  and g22896 (n12173, n11862, n12171);
  not g22897 (n_10982, n12172);
  not g22898 (n_10983, n12173);
  and g22899 (n12174, n_10982, n_10983);
  not g22900 (n_10984, n12159);
  and g22901 (n12175, n_10984, n12174);
  not g22902 (n_10985, n12175);
  and g22903 (n12176, n_10984, n_10985);
  and g22904 (n12177, n12174, n_10985);
  not g22905 (n_10986, n12176);
  not g22906 (n_10987, n12177);
  and g22907 (n12178, n_10986, n_10987);
  not g22908 (n_10988, n12146);
  not g22909 (n_10989, n12178);
  and g22910 (n12179, n_10988, n_10989);
  not g22911 (n_10990, n12179);
  and g22912 (n12180, n_10988, n_10990);
  and g22913 (n12181, n_10989, n_10990);
  not g22914 (n_10991, n12180);
  not g22915 (n_10992, n12181);
  and g22916 (n12182, n_10991, n_10992);
  and g22917 (n12183, n_10655, n_10659);
  and g22918 (n12184, n12182, n12183);
  not g22919 (n_10993, n12182);
  not g22920 (n_10994, n12183);
  and g22921 (n12185, n_10993, n_10994);
  not g22922 (n_10995, n12184);
  not g22923 (n_10996, n12185);
  and g22924 (n12186, n_10995, n_10996);
  and g22925 (n12187, n_10634, n_10639);
  and g22926 (n12188, n11953, n11968);
  not g22927 (n_10997, n11953);
  not g22928 (n_10998, n11968);
  and g22929 (n12189, n_10997, n_10998);
  not g22930 (n_10999, n12188);
  not g22931 (n_11000, n12189);
  and g22932 (n12190, n_10999, n_11000);
  not g22933 (n_11001, n12190);
  and g22934 (n12191, n11785, n_11001);
  not g22935 (n_11002, n11785);
  and g22936 (n12192, n_11002, n12190);
  not g22937 (n_11003, n12191);
  not g22938 (n_11004, n12192);
  and g22939 (n12193, n_11003, n_11004);
  and g22940 (n12194, n_10625, n_10631);
  not g22941 (n_11005, n12193);
  and g22942 (n12195, n_11005, n12194);
  not g22943 (n_11006, n12194);
  and g22944 (n12196, n12193, n_11006);
  not g22945 (n_11007, n12195);
  not g22946 (n_11008, n12196);
  and g22947 (n12197, n_11007, n_11008);
  and g22948 (n12198, \a[10] , \a[63] );
  and g22949 (n12199, \a[12] , \a[61] );
  not g22950 (n_11009, n12198);
  not g22951 (n_11010, n12199);
  and g22952 (n12200, n_11009, n_11010);
  and g22953 (n12201, n480, n9909);
  not g22954 (n_11011, n12201);
  not g22957 (n_11012, n12200);
  not g22959 (n_11013, n12204);
  and g22960 (n12205, n_11011, n_11013);
  and g22961 (n12206, n_11012, n12205);
  and g22962 (n12207, \a[48] , n_11013);
  and g22963 (n12208, \a[25] , n12207);
  not g22964 (n_11014, n12206);
  not g22965 (n_11015, n12208);
  and g22966 (n12209, n_11014, n_11015);
  and g22967 (n12210, n2617, n5296);
  and g22968 (n12211, n3110, n4811);
  and g22969 (n12212, n2334, n5713);
  not g22970 (n_11016, n12211);
  not g22971 (n_11017, n12212);
  and g22972 (n12213, n_11016, n_11017);
  not g22973 (n_11018, n12210);
  not g22974 (n_11019, n12213);
  and g22975 (n12214, n_11018, n_11019);
  not g22976 (n_11020, n12214);
  and g22977 (n12215, \a[45] , n_11020);
  and g22978 (n12216, \a[28] , n12215);
  and g22979 (n12217, n_11018, n_11020);
  and g22980 (n12218, \a[29] , \a[44] );
  and g22981 (n12219, \a[30] , \a[43] );
  not g22982 (n_11021, n12218);
  not g22983 (n_11022, n12219);
  and g22984 (n12220, n_11021, n_11022);
  not g22985 (n_11023, n12220);
  and g22986 (n12221, n12217, n_11023);
  not g22987 (n_11024, n12216);
  not g22988 (n_11025, n12221);
  and g22989 (n12222, n_11024, n_11025);
  not g22990 (n_11026, n12209);
  not g22991 (n_11027, n12222);
  and g22992 (n12223, n_11026, n_11027);
  not g22993 (n_11028, n12223);
  and g22994 (n12224, n_11026, n_11028);
  and g22995 (n12225, n_11027, n_11028);
  not g22996 (n_11029, n12224);
  not g22997 (n_11030, n12225);
  and g22998 (n12226, n_11029, n_11030);
  and g22999 (n12227, n3828, n4565);
  and g23000 (n12228, n3687, n4748);
  and g23001 (n12229, n3319, n5083);
  not g23002 (n_11031, n12228);
  not g23003 (n_11032, n12229);
  and g23004 (n12230, n_11031, n_11032);
  not g23005 (n_11033, n12227);
  not g23006 (n_11034, n12230);
  and g23007 (n12231, n_11033, n_11034);
  not g23008 (n_11035, n12231);
  and g23009 (n12232, n4748, n_11035);
  and g23010 (n12233, n_11033, n_11035);
  and g23011 (n12234, \a[35] , \a[38] );
  not g23012 (n_11036, n3687);
  not g23013 (n_11037, n12234);
  and g23014 (n12235, n_11036, n_11037);
  not g23015 (n_11038, n12235);
  and g23016 (n12236, n12233, n_11038);
  not g23017 (n_11039, n12232);
  not g23018 (n_11040, n12236);
  and g23019 (n12237, n_11039, n_11040);
  not g23020 (n_11041, n12226);
  not g23021 (n_11042, n12237);
  and g23022 (n12238, n_11041, n_11042);
  not g23023 (n_11043, n12238);
  and g23024 (n12239, n_11041, n_11043);
  and g23025 (n12240, n_11042, n_11043);
  not g23026 (n_11044, n12239);
  not g23027 (n_11045, n12240);
  and g23028 (n12241, n_11044, n_11045);
  not g23029 (n_11046, n12197);
  and g23030 (n12242, n_11046, n12241);
  not g23031 (n_11047, n12241);
  and g23032 (n12243, n12197, n_11047);
  not g23033 (n_11048, n12242);
  not g23034 (n_11049, n12243);
  and g23035 (n12244, n_11048, n_11049);
  not g23036 (n_11050, n12187);
  and g23037 (n12245, n_11050, n12244);
  not g23038 (n_11051, n12245);
  and g23039 (n12246, n_11050, n_11051);
  and g23040 (n12247, n12244, n_11051);
  not g23041 (n_11052, n12246);
  not g23042 (n_11053, n12247);
  and g23043 (n12248, n_11052, n_11053);
  not g23044 (n_11054, n12248);
  and g23045 (n12249, n12186, n_11054);
  not g23046 (n_11055, n12249);
  and g23047 (n12250, n12186, n_11055);
  and g23048 (n12251, n_11054, n_11055);
  not g23049 (n_11056, n12250);
  not g23050 (n_11057, n12251);
  and g23051 (n12252, n_11056, n_11057);
  not g23052 (n_11058, n12252);
  and g23053 (n12253, n12101, n_11058);
  not g23054 (n_11059, n12253);
  and g23055 (n12254, n12101, n_11059);
  and g23056 (n12255, n_11058, n_11059);
  not g23057 (n_11060, n12254);
  not g23058 (n_11061, n12255);
  and g23059 (n12256, n_11060, n_11061);
  not g23060 (n_11062, n12061);
  and g23061 (n12257, n_11062, n12256);
  not g23062 (n_11063, n12256);
  and g23063 (n12258, n12061, n_11063);
  not g23064 (n_11064, n12257);
  not g23065 (n_11065, n12258);
  and g23066 (n12259, n_11064, n_11065);
  not g23067 (n_11066, n12259);
  and g23068 (n12260, n12019, n_11066);
  not g23069 (n_11067, n12019);
  and g23070 (n12261, n_11067, n12259);
  not g23071 (n_11068, n12260);
  not g23072 (n_11069, n12261);
  and g23073 (n12262, n_11068, n_11069);
  not g23074 (n_11070, n12018);
  not g23075 (n_11071, n12262);
  and g23076 (n12263, n_11070, n_11071);
  and g23077 (n12264, n12018, n12262);
  or g23078 (\asquared[74] , n12263, n12264);
  and g23079 (n12266, n_10881, n_11065);
  and g23080 (n12267, n_10872, n_10876);
  and g23081 (n12268, n12032, n12233);
  not g23082 (n_11072, n12032);
  not g23083 (n_11073, n12233);
  and g23084 (n12269, n_11072, n_11073);
  not g23085 (n_11074, n12268);
  not g23086 (n_11075, n12269);
  and g23087 (n12270, n_11074, n_11075);
  and g23088 (n12271, n891, n8987);
  and g23089 (n12272, n893, n10089);
  and g23090 (n12273, n895, n9509);
  not g23091 (n_11076, n12272);
  not g23092 (n_11077, n12273);
  and g23093 (n12274, n_11076, n_11077);
  not g23094 (n_11078, n12271);
  not g23095 (n_11079, n12274);
  and g23096 (n12275, n_11078, n_11079);
  not g23097 (n_11080, n12275);
  and g23098 (n12276, \a[60] , n_11080);
  and g23099 (n12277, \a[14] , n12276);
  and g23100 (n12278, \a[15] , \a[59] );
  and g23101 (n12279, \a[16] , \a[58] );
  not g23102 (n_11081, n12278);
  not g23103 (n_11082, n12279);
  and g23104 (n12280, n_11081, n_11082);
  and g23105 (n12281, n_11078, n_11080);
  not g23106 (n_11083, n12280);
  and g23107 (n12282, n_11083, n12281);
  not g23108 (n_11084, n12277);
  not g23109 (n_11085, n12282);
  and g23110 (n12283, n_11084, n_11085);
  not g23111 (n_11086, n12283);
  and g23112 (n12284, n12270, n_11086);
  not g23113 (n_11087, n12284);
  and g23114 (n12285, n12270, n_11087);
  and g23115 (n12286, n_11086, n_11087);
  not g23116 (n_11088, n12285);
  not g23117 (n_11089, n12286);
  and g23118 (n12287, n_11088, n_11089);
  and g23119 (n12288, n_10945, n_10960);
  and g23120 (n12289, n12287, n12288);
  not g23121 (n_11090, n12287);
  not g23122 (n_11091, n12288);
  and g23123 (n12290, n_11090, n_11091);
  not g23124 (n_11092, n12289);
  not g23125 (n_11093, n12290);
  and g23126 (n12291, n_11092, n_11093);
  and g23127 (n12292, n_10855, n_10861);
  not g23128 (n_11094, n12291);
  and g23129 (n12293, n_11094, n12292);
  not g23130 (n_11095, n12292);
  and g23131 (n12294, n12291, n_11095);
  not g23132 (n_11096, n12293);
  not g23133 (n_11097, n12294);
  and g23134 (n12295, n_11096, n_11097);
  and g23135 (n12296, n_10990, n_10996);
  and g23136 (n12297, n_11008, n_11049);
  not g23137 (n_11098, n12296);
  not g23138 (n_11099, n12297);
  and g23139 (n12298, n_11098, n_11099);
  not g23140 (n_11100, n12298);
  and g23141 (n12299, n_11098, n_11100);
  and g23142 (n12300, n_11099, n_11100);
  not g23143 (n_11101, n12299);
  not g23144 (n_11102, n12300);
  and g23145 (n12301, n_11101, n_11102);
  not g23146 (n_11103, n12301);
  and g23147 (n12302, n12295, n_11103);
  not g23148 (n_11104, n12295);
  and g23149 (n12303, n_11104, n12301);
  not g23150 (n_11105, n12267);
  not g23151 (n_11106, n12303);
  and g23152 (n12304, n_11105, n_11106);
  not g23153 (n_11107, n12302);
  and g23154 (n12305, n_11107, n12304);
  not g23155 (n_11108, n12305);
  and g23156 (n12306, n_11105, n_11108);
  and g23157 (n12307, n_11106, n_11108);
  and g23158 (n12308, n_11107, n12307);
  not g23159 (n_11109, n12306);
  not g23160 (n_11110, n12308);
  and g23161 (n12309, n_11109, n_11110);
  and g23162 (n12310, n748, n9721);
  not g23163 (n_11111, n12310);
  and g23164 (n12311, \a[61] , n_11111);
  and g23165 (n12312, \a[13] , n12311);
  and g23166 (n12313, \a[62] , n_11111);
  and g23167 (n12314, \a[12] , n12313);
  not g23168 (n_11112, n12312);
  not g23169 (n_11113, n12314);
  and g23170 (n12315, n_11112, n_11113);
  not g23171 (n_11114, n12108);
  not g23172 (n_11115, n12315);
  and g23173 (n12316, n_11114, n_11115);
  not g23174 (n_11116, n12316);
  and g23175 (n12317, n_11114, n_11116);
  and g23176 (n12318, n_11115, n_11116);
  not g23177 (n_11117, n12317);
  not g23178 (n_11118, n12318);
  and g23179 (n12319, n_11117, n_11118);
  and g23180 (n12320, \a[30] , \a[44] );
  and g23181 (n12321, n9618, n12320);
  and g23182 (n12322, n2617, n5713);
  and g23183 (n12323, \a[29] , \a[57] );
  and g23184 (n12324, n9119, n12323);
  not g23185 (n_11119, n12322);
  not g23186 (n_11120, n12324);
  and g23187 (n12325, n_11119, n_11120);
  not g23188 (n_11121, n12321);
  not g23189 (n_11122, n12325);
  and g23190 (n12326, n_11121, n_11122);
  not g23191 (n_11123, n12326);
  and g23192 (n12327, \a[45] , n_11123);
  and g23193 (n12328, \a[29] , n12327);
  and g23194 (n12329, n_11121, n_11123);
  not g23195 (n_11124, n9618);
  not g23196 (n_11125, n12320);
  and g23197 (n12330, n_11124, n_11125);
  not g23198 (n_11126, n12330);
  and g23199 (n12331, n12329, n_11126);
  not g23200 (n_11127, n12328);
  not g23201 (n_11128, n12331);
  and g23202 (n12332, n_11127, n_11128);
  not g23203 (n_11129, n12319);
  not g23204 (n_11130, n12332);
  and g23205 (n12333, n_11129, n_11130);
  not g23206 (n_11131, n12333);
  and g23207 (n12334, n_11129, n_11131);
  and g23208 (n12335, n_11130, n_11131);
  not g23209 (n_11132, n12334);
  not g23210 (n_11133, n12335);
  and g23211 (n12336, n_11132, n_11133);
  and g23212 (n12337, n_11000, n_11004);
  and g23213 (n12338, n12336, n12337);
  not g23214 (n_11134, n12336);
  not g23215 (n_11135, n12337);
  and g23216 (n12339, n_11134, n_11135);
  not g23217 (n_11136, n12338);
  not g23218 (n_11137, n12339);
  and g23219 (n12340, n_11136, n_11137);
  and g23220 (n12341, \a[31] , \a[43] );
  and g23221 (n12342, \a[32] , \a[42] );
  not g23222 (n_11138, n12341);
  not g23223 (n_11139, n12342);
  and g23224 (n12343, n_11138, n_11139);
  and g23225 (n12344, n3812, n5018);
  not g23226 (n_11140, n12344);
  not g23228 (n_11141, n12343);
  not g23231 (n_11142, n12347);
  and g23232 (n12348, n_11140, n_11142);
  and g23233 (n12349, n_11141, n12348);
  and g23234 (n12350, \a[63] , n_11142);
  and g23235 (n12351, \a[11] , n12350);
  not g23236 (n_11143, n12349);
  not g23237 (n_11144, n12351);
  and g23238 (n12352, n_11143, n_11144);
  and g23239 (n12353, \a[18] , \a[56] );
  and g23240 (n12354, \a[25] , \a[49] );
  not g23241 (n_11145, n12353);
  not g23242 (n_11146, n12354);
  and g23243 (n12355, n_11145, n_11146);
  and g23244 (n12356, \a[25] , \a[56] );
  and g23245 (n12357, n10490, n12356);
  not g23246 (n_11147, n12357);
  and g23247 (n12358, n5342, n_11147);
  not g23248 (n_11148, n12355);
  and g23249 (n12359, n_11148, n12358);
  not g23250 (n_11149, n12359);
  and g23251 (n12360, n5342, n_11149);
  and g23252 (n12361, n_11147, n_11149);
  and g23253 (n12362, n_11148, n12361);
  not g23254 (n_11150, n12360);
  not g23255 (n_11151, n12362);
  and g23256 (n12363, n_11150, n_11151);
  not g23257 (n_11152, n12352);
  not g23258 (n_11153, n12363);
  and g23259 (n12364, n_11152, n_11153);
  not g23260 (n_11154, n12364);
  and g23261 (n12365, n_11152, n_11154);
  and g23262 (n12366, n_11153, n_11154);
  not g23263 (n_11155, n12365);
  not g23264 (n_11156, n12366);
  and g23265 (n12367, n_11155, n_11156);
  and g23266 (n12368, n2331, n5666);
  and g23267 (n12369, n2800, n8578);
  and g23268 (n12370, n2227, n6252);
  not g23269 (n_11157, n12369);
  not g23270 (n_11158, n12370);
  and g23271 (n12371, n_11157, n_11158);
  not g23272 (n_11159, n12368);
  not g23273 (n_11160, n12371);
  and g23274 (n12372, n_11159, n_11160);
  not g23275 (n_11161, n12372);
  and g23276 (n12373, \a[48] , n_11161);
  and g23277 (n12374, \a[26] , n12373);
  and g23278 (n12375, n_11159, n_11161);
  and g23279 (n12376, \a[27] , \a[47] );
  and g23280 (n12377, \a[28] , \a[46] );
  not g23281 (n_11162, n12376);
  not g23282 (n_11163, n12377);
  and g23283 (n12378, n_11162, n_11163);
  not g23284 (n_11164, n12378);
  and g23285 (n12379, n12375, n_11164);
  not g23286 (n_11165, n12374);
  not g23287 (n_11166, n12379);
  and g23288 (n12380, n_11165, n_11166);
  not g23289 (n_11167, n12367);
  not g23290 (n_11168, n12380);
  and g23291 (n12381, n_11167, n_11168);
  not g23292 (n_11169, n12381);
  and g23293 (n12382, n_11167, n_11169);
  and g23294 (n12383, n_11168, n_11169);
  not g23295 (n_11170, n12382);
  not g23296 (n_11171, n12383);
  and g23297 (n12384, n_11170, n_11171);
  and g23298 (n12385, \a[21] , \a[53] );
  not g23299 (n_11172, n8212);
  not g23300 (n_11173, n12385);
  and g23301 (n12386, n_11172, n_11173);
  and g23302 (n12387, n1492, n7697);
  and g23303 (n12388, \a[52] , \a[55] );
  and g23304 (n12389, n4036, n12388);
  and g23305 (n12390, n1574, n7433);
  not g23306 (n_11174, n12389);
  not g23307 (n_11175, n12390);
  and g23308 (n12391, n_11174, n_11175);
  not g23309 (n_11176, n12387);
  not g23310 (n_11177, n12391);
  and g23311 (n12392, n_11176, n_11177);
  not g23312 (n_11178, n12392);
  and g23313 (n12393, n_11176, n_11178);
  not g23314 (n_11179, n12386);
  and g23315 (n12394, n_11179, n12393);
  and g23316 (n12395, \a[52] , n_11178);
  and g23317 (n12396, \a[22] , n12395);
  not g23318 (n_11180, n12394);
  not g23319 (n_11181, n12396);
  and g23320 (n12397, n_11180, n_11181);
  and g23321 (n12398, \a[35] , \a[39] );
  not g23322 (n_11182, n5195);
  not g23323 (n_11183, n12398);
  and g23324 (n12399, n_11182, n_11183);
  and g23325 (n12400, n3319, n4171);
  not g23326 (n_11184, n12400);
  and g23327 (n12401, n11043, n_11184);
  not g23328 (n_11185, n12399);
  and g23329 (n12402, n_11185, n12401);
  not g23330 (n_11186, n12402);
  and g23331 (n12403, n11043, n_11186);
  and g23332 (n12404, n_11184, n_11186);
  and g23333 (n12405, n_11185, n12404);
  not g23334 (n_11187, n12403);
  not g23335 (n_11188, n12405);
  and g23336 (n12406, n_11187, n_11188);
  not g23337 (n_11189, n12397);
  not g23338 (n_11190, n12406);
  and g23339 (n12407, n_11189, n_11190);
  not g23340 (n_11191, n12407);
  and g23341 (n12408, n_11189, n_11191);
  and g23342 (n12409, n_11190, n_11191);
  not g23343 (n_11192, n12408);
  not g23344 (n_11193, n12409);
  and g23345 (n12410, n_11192, n_11193);
  and g23346 (n12411, \a[23] , \a[51] );
  and g23347 (n12412, \a[24] , \a[50] );
  not g23348 (n_11194, n12411);
  not g23349 (n_11195, n12412);
  and g23350 (n12413, n_11194, n_11195);
  and g23351 (n12414, n1666, n6564);
  not g23352 (n_11196, n12414);
  and g23353 (n12415, n3530, n_11196);
  not g23354 (n_11197, n12413);
  and g23355 (n12416, n_11197, n12415);
  not g23356 (n_11198, n12416);
  and g23357 (n12417, n3530, n_11198);
  and g23358 (n12418, n_11196, n_11198);
  and g23359 (n12419, n_11197, n12418);
  not g23360 (n_11199, n12417);
  not g23361 (n_11200, n12419);
  and g23362 (n12420, n_11199, n_11200);
  not g23363 (n_11201, n12410);
  not g23364 (n_11202, n12420);
  and g23365 (n12421, n_11201, n_11202);
  not g23366 (n_11203, n12421);
  and g23367 (n12422, n_11201, n_11203);
  and g23368 (n12423, n_11202, n_11203);
  not g23369 (n_11204, n12422);
  not g23370 (n_11205, n12423);
  and g23371 (n12424, n_11204, n_11205);
  not g23372 (n_11206, n12384);
  and g23373 (n12425, n_11206, n12424);
  not g23374 (n_11207, n12424);
  and g23375 (n12426, n12384, n_11207);
  not g23376 (n_11208, n12425);
  not g23377 (n_11209, n12426);
  and g23378 (n12427, n_11208, n_11209);
  not g23379 (n_11210, n12427);
  and g23380 (n12428, n12340, n_11210);
  not g23381 (n_11211, n12428);
  and g23382 (n12429, n12340, n_11211);
  and g23383 (n12430, n_11210, n_11211);
  not g23384 (n_11212, n12429);
  not g23385 (n_11213, n12430);
  and g23386 (n12431, n_11212, n_11213);
  and g23387 (n12432, n_10864, n_10868);
  and g23388 (n12433, n12169, n12217);
  not g23389 (n_11214, n12169);
  not g23390 (n_11215, n12217);
  and g23391 (n12434, n_11214, n_11215);
  not g23392 (n_11216, n12433);
  not g23393 (n_11217, n12434);
  and g23394 (n12435, n_11216, n_11217);
  not g23395 (n_11218, n12435);
  and g23396 (n12436, n12155, n_11218);
  not g23397 (n_11219, n12155);
  and g23398 (n12437, n_11219, n12435);
  not g23399 (n_11220, n12436);
  not g23400 (n_11221, n12437);
  and g23401 (n12438, n_11220, n_11221);
  and g23402 (n12439, n12121, n12137);
  not g23403 (n_11222, n12121);
  not g23404 (n_11223, n12137);
  and g23405 (n12440, n_11222, n_11223);
  not g23406 (n_11224, n12439);
  not g23407 (n_11225, n12440);
  and g23408 (n12441, n_11224, n_11225);
  not g23409 (n_11226, n12441);
  and g23410 (n12442, n12205, n_11226);
  not g23411 (n_11227, n12205);
  and g23412 (n12443, n_11227, n12441);
  not g23413 (n_11228, n12442);
  not g23414 (n_11229, n12443);
  and g23415 (n12444, n_11228, n_11229);
  and g23416 (n12445, n_11028, n_11043);
  not g23417 (n_11230, n12444);
  and g23418 (n12446, n_11230, n12445);
  not g23419 (n_11231, n12445);
  and g23420 (n12447, n12444, n_11231);
  not g23421 (n_11232, n12446);
  not g23422 (n_11233, n12447);
  and g23423 (n12448, n_11232, n_11233);
  and g23424 (n12449, n12438, n12448);
  not g23425 (n_11234, n12438);
  not g23426 (n_11235, n12448);
  and g23427 (n12450, n_11234, n_11235);
  not g23428 (n_11236, n12449);
  not g23429 (n_11237, n12450);
  and g23430 (n12451, n_11236, n_11237);
  not g23431 (n_11238, n12432);
  and g23432 (n12452, n_11238, n12451);
  not g23433 (n_11239, n12451);
  and g23434 (n12453, n12432, n_11239);
  not g23435 (n_11240, n12452);
  not g23436 (n_11241, n12453);
  and g23437 (n12454, n_11240, n_11241);
  not g23438 (n_11242, n12431);
  and g23439 (n12455, n_11242, n12454);
  not g23440 (n_11243, n12455);
  and g23441 (n12456, n12454, n_11243);
  and g23442 (n12457, n_11242, n_11243);
  not g23443 (n_11244, n12456);
  not g23444 (n_11245, n12457);
  and g23445 (n12458, n_11244, n_11245);
  not g23446 (n_11246, n12309);
  and g23447 (n12459, n_11246, n12458);
  not g23448 (n_11247, n12458);
  and g23449 (n12460, n12309, n_11247);
  not g23450 (n_11248, n12459);
  not g23451 (n_11249, n12460);
  and g23452 (n12461, n_11248, n_11249);
  and g23453 (n12462, n_10925, n_11059);
  and g23454 (n12463, n_11051, n_11055);
  and g23455 (n12464, n_10893, n_10920);
  and g23456 (n12465, n_10905, n_10909);
  and g23457 (n12466, n_10896, n_10901);
  and g23458 (n12467, n12465, n12466);
  not g23459 (n_11250, n12465);
  not g23460 (n_11251, n12466);
  and g23461 (n12468, n_11250, n_11251);
  not g23462 (n_11252, n12467);
  not g23463 (n_11253, n12468);
  and g23464 (n12469, n_11252, n_11253);
  and g23465 (n12470, n_10982, n_10985);
  not g23466 (n_11254, n12469);
  and g23467 (n12471, n_11254, n12470);
  not g23468 (n_11255, n12470);
  and g23469 (n12472, n12469, n_11255);
  not g23470 (n_11256, n12471);
  not g23471 (n_11257, n12472);
  and g23472 (n12473, n_11256, n_11257);
  and g23473 (n12474, n_10912, n_10916);
  and g23474 (n12475, n_10885, n_10889);
  and g23475 (n12476, n12474, n12475);
  not g23476 (n_11258, n12474);
  not g23477 (n_11259, n12475);
  and g23478 (n12477, n_11258, n_11259);
  not g23479 (n_11260, n12476);
  not g23480 (n_11261, n12477);
  and g23481 (n12478, n_11260, n_11261);
  and g23482 (n12479, n12473, n12478);
  not g23483 (n_11262, n12473);
  not g23484 (n_11263, n12478);
  and g23485 (n12480, n_11262, n_11263);
  not g23486 (n_11264, n12479);
  not g23487 (n_11265, n12480);
  and g23488 (n12481, n_11264, n_11265);
  not g23489 (n_11266, n12464);
  and g23490 (n12482, n_11266, n12481);
  not g23491 (n_11267, n12481);
  and g23492 (n12483, n12464, n_11267);
  not g23493 (n_11268, n12482);
  not g23494 (n_11269, n12483);
  and g23495 (n12484, n_11268, n_11269);
  not g23496 (n_11270, n12463);
  and g23497 (n12485, n_11270, n12484);
  not g23498 (n_11271, n12484);
  and g23499 (n12486, n12463, n_11271);
  not g23500 (n_11272, n12485);
  not g23501 (n_11273, n12486);
  and g23502 (n12487, n_11272, n_11273);
  not g23503 (n_11274, n12462);
  and g23504 (n12488, n_11274, n12487);
  not g23505 (n_11275, n12487);
  and g23506 (n12489, n12462, n_11275);
  not g23507 (n_11276, n12488);
  not g23508 (n_11277, n12489);
  and g23509 (n12490, n_11276, n_11277);
  not g23510 (n_11278, n12461);
  and g23511 (n12491, n_11278, n12490);
  not g23512 (n_11279, n12490);
  and g23513 (n12492, n12461, n_11279);
  not g23514 (n_11280, n12491);
  not g23515 (n_11281, n12492);
  and g23516 (n12493, n_11280, n_11281);
  not g23517 (n_11282, n12493);
  and g23518 (n12494, n12266, n_11282);
  not g23519 (n_11283, n12266);
  and g23520 (n12495, n_11283, n12493);
  not g23521 (n_11284, n12494);
  not g23522 (n_11285, n12495);
  and g23523 (n12496, n_11284, n_11285);
  and g23524 (n12497, n_11070, n_11068);
  not g23525 (n_11286, n12497);
  and g23526 (n12498, n_11069, n_11286);
  not g23527 (n_11287, n12496);
  and g23528 (n12499, n_11287, n12498);
  not g23529 (n_11288, n12498);
  and g23530 (n12500, n12496, n_11288);
  not g23531 (n_11289, n12499);
  not g23532 (n_11290, n12500);
  and g23533 (\asquared[75] , n_11289, n_11290);
  and g23534 (n12502, n_11276, n_11280);
  and g23535 (n12503, n_11268, n_11272);
  and g23536 (n12504, n_11075, n_11087);
  and g23537 (n12505, n_11225, n_11229);
  and g23538 (n12506, n12504, n12505);
  not g23539 (n_11291, n12504);
  not g23540 (n_11292, n12505);
  and g23541 (n12507, n_11291, n_11292);
  not g23542 (n_11293, n12506);
  not g23543 (n_11294, n12507);
  and g23544 (n12508, n_11293, n_11294);
  and g23545 (n12509, n_11217, n_11221);
  not g23546 (n_11295, n12508);
  and g23547 (n12510, n_11295, n12509);
  not g23548 (n_11296, n12509);
  and g23549 (n12511, n12508, n_11296);
  not g23550 (n_11297, n12510);
  not g23551 (n_11298, n12511);
  and g23552 (n12512, n_11297, n_11298);
  and g23553 (n12513, n_11206, n_11207);
  not g23554 (n_11299, n12513);
  and g23555 (n12514, n_11211, n_11299);
  not g23556 (n_11300, n12514);
  and g23557 (n12515, n12512, n_11300);
  not g23558 (n_11301, n12512);
  and g23559 (n12516, n_11301, n12514);
  not g23560 (n_11302, n12515);
  not g23561 (n_11303, n12516);
  and g23562 (n12517, n_11302, n_11303);
  and g23563 (n12518, n_11131, n_11137);
  and g23564 (n12519, n12404, n12418);
  not g23565 (n_11304, n12404);
  not g23566 (n_11305, n12418);
  and g23567 (n12520, n_11304, n_11305);
  not g23568 (n_11306, n12519);
  not g23569 (n_11307, n12520);
  and g23570 (n12521, n_11306, n_11307);
  not g23571 (n_11308, n12521);
  and g23572 (n12522, n12393, n_11308);
  not g23573 (n_11309, n12393);
  and g23574 (n12523, n_11309, n12521);
  not g23575 (n_11310, n12522);
  not g23576 (n_11311, n12523);
  and g23577 (n12524, n_11310, n_11311);
  and g23578 (n12525, n12348, n12361);
  not g23579 (n_11312, n12348);
  not g23580 (n_11313, n12361);
  and g23581 (n12526, n_11312, n_11313);
  not g23582 (n_11314, n12525);
  not g23583 (n_11315, n12526);
  and g23584 (n12527, n_11314, n_11315);
  and g23585 (n12528, n_11111, n_11116);
  not g23586 (n_11316, n12527);
  and g23587 (n12529, n_11316, n12528);
  not g23588 (n_11317, n12528);
  and g23589 (n12530, n12527, n_11317);
  not g23590 (n_11318, n12529);
  not g23591 (n_11319, n12530);
  and g23592 (n12531, n_11318, n_11319);
  and g23593 (n12532, n12524, n12531);
  not g23594 (n_11320, n12524);
  not g23595 (n_11321, n12531);
  and g23596 (n12533, n_11320, n_11321);
  not g23597 (n_11322, n12532);
  not g23598 (n_11323, n12533);
  and g23599 (n12534, n_11322, n_11323);
  not g23600 (n_11324, n12518);
  and g23601 (n12535, n_11324, n12534);
  not g23602 (n_11325, n12534);
  and g23603 (n12536, n12518, n_11325);
  not g23604 (n_11326, n12535);
  not g23605 (n_11327, n12536);
  and g23606 (n12537, n_11326, n_11327);
  and g23607 (n12538, n12517, n12537);
  not g23608 (n_11328, n12517);
  not g23609 (n_11329, n12537);
  and g23610 (n12539, n_11328, n_11329);
  not g23611 (n_11330, n12538);
  not g23612 (n_11331, n12539);
  and g23613 (n12540, n_11330, n_11331);
  not g23614 (n_11332, n12540);
  and g23615 (n12541, n12503, n_11332);
  not g23616 (n_11333, n12503);
  and g23617 (n12542, n_11333, n12540);
  not g23618 (n_11334, n12541);
  not g23619 (n_11335, n12542);
  and g23620 (n12543, n_11334, n_11335);
  and g23621 (n12544, \a[12] , \a[63] );
  and g23622 (n12545, \a[19] , \a[56] );
  not g23623 (n_11336, n12544);
  not g23624 (n_11337, n12545);
  and g23625 (n12546, n_11336, n_11337);
  and g23626 (n12547, \a[19] , \a[63] );
  and g23627 (n12548, n10885, n12547);
  not g23628 (n_11338, n12548);
  not g23631 (n_11339, n12546);
  not g23633 (n_11340, n12551);
  and g23634 (n12552, n_11338, n_11340);
  and g23635 (n12553, n_11339, n12552);
  and g23636 (n12554, \a[45] , n_11340);
  and g23637 (n12555, \a[30] , n12554);
  not g23638 (n_11341, n12553);
  not g23639 (n_11342, n12555);
  and g23640 (n12556, n_11341, n_11342);
  and g23641 (n12557, \a[23] , \a[52] );
  and g23642 (n12558, \a[35] , \a[40] );
  not g23643 (n_11343, n8936);
  not g23644 (n_11344, n12558);
  and g23645 (n12559, n_11343, n_11344);
  and g23646 (n12560, n3828, n4171);
  not g23647 (n_11345, n12560);
  and g23648 (n12561, n12557, n_11345);
  not g23649 (n_11346, n12559);
  and g23650 (n12562, n_11346, n12561);
  not g23651 (n_11347, n12562);
  and g23652 (n12563, n12557, n_11347);
  and g23653 (n12564, n_11345, n_11347);
  and g23654 (n12565, n_11346, n12564);
  not g23655 (n_11348, n12563);
  not g23656 (n_11349, n12565);
  and g23657 (n12566, n_11348, n_11349);
  not g23658 (n_11350, n12556);
  not g23659 (n_11351, n12566);
  and g23660 (n12567, n_11350, n_11351);
  not g23661 (n_11352, n12567);
  and g23662 (n12568, n_11350, n_11352);
  and g23663 (n12569, n_11351, n_11352);
  not g23664 (n_11353, n12568);
  not g23665 (n_11354, n12569);
  and g23666 (n12570, n_11353, n_11354);
  and g23667 (n12571, \a[38] , \a[62] );
  and g23668 (n12572, \a[13] , n12571);
  not g23669 (n_11355, n12572);
  and g23670 (n12573, n4565, n_11355);
  not g23671 (n_11356, n12573);
  and g23672 (n12574, n4565, n_11356);
  and g23673 (n12575, n_11355, n_11356);
  and g23674 (n12576, \a[13] , \a[62] );
  not g23675 (n_11357, \a[38] );
  not g23676 (n_11358, n12576);
  and g23677 (n12577, n_11357, n_11358);
  not g23678 (n_11359, n12577);
  and g23679 (n12578, n12575, n_11359);
  not g23680 (n_11360, n12574);
  not g23681 (n_11361, n12578);
  and g23682 (n12579, n_11360, n_11361);
  not g23683 (n_11362, n12570);
  not g23684 (n_11363, n12579);
  and g23685 (n12580, n_11362, n_11363);
  not g23686 (n_11364, n12580);
  and g23687 (n12581, n_11362, n_11364);
  and g23688 (n12582, n_11363, n_11364);
  not g23689 (n_11365, n12581);
  not g23690 (n_11366, n12582);
  and g23691 (n12583, n_11365, n_11366);
  and g23692 (n12584, n_11253, n_11257);
  and g23693 (n12585, n12583, n12584);
  not g23694 (n_11367, n12583);
  not g23695 (n_11368, n12584);
  and g23696 (n12586, n_11367, n_11368);
  not g23697 (n_11369, n12585);
  not g23698 (n_11370, n12586);
  and g23699 (n12587, n_11369, n_11370);
  and g23700 (n12588, n891, n9509);
  and g23701 (n12589, n893, n8905);
  and g23702 (n12590, n895, n9512);
  not g23703 (n_11371, n12589);
  not g23704 (n_11372, n12590);
  and g23705 (n12591, n_11371, n_11372);
  not g23706 (n_11373, n12588);
  not g23707 (n_11374, n12591);
  and g23708 (n12592, n_11373, n_11374);
  not g23709 (n_11375, n12592);
  and g23710 (n12593, n_11373, n_11375);
  and g23711 (n12594, \a[15] , \a[60] );
  and g23712 (n12595, \a[16] , \a[59] );
  not g23713 (n_11376, n12594);
  not g23714 (n_11377, n12595);
  and g23715 (n12596, n_11376, n_11377);
  not g23716 (n_11378, n12596);
  and g23717 (n12597, n12593, n_11378);
  and g23718 (n12598, \a[61] , n_11375);
  and g23719 (n12599, \a[14] , n12598);
  not g23720 (n_11379, n12597);
  not g23721 (n_11380, n12599);
  and g23722 (n12600, n_11379, n_11380);
  and g23723 (n12601, \a[49] , \a[57] );
  and g23724 (n12602, n4543, n12601);
  and g23725 (n12603, \a[26] , \a[58] );
  and g23726 (n12604, n7063, n12603);
  and g23727 (n12605, n1052, n8436);
  not g23728 (n_11381, n12604);
  not g23729 (n_11382, n12605);
  and g23730 (n12606, n_11381, n_11382);
  not g23731 (n_11383, n12602);
  not g23732 (n_11384, n12606);
  and g23733 (n12607, n_11383, n_11384);
  not g23734 (n_11385, n12607);
  and g23735 (n12608, \a[58] , n_11385);
  and g23736 (n12609, \a[17] , n12608);
  and g23737 (n12610, n_11383, n_11385);
  and g23738 (n12611, \a[18] , \a[57] );
  and g23739 (n12612, \a[26] , \a[49] );
  not g23740 (n_11386, n12611);
  not g23741 (n_11387, n12612);
  and g23742 (n12613, n_11386, n_11387);
  not g23743 (n_11388, n12613);
  and g23744 (n12614, n12610, n_11388);
  not g23745 (n_11389, n12609);
  not g23746 (n_11390, n12614);
  and g23747 (n12615, n_11389, n_11390);
  not g23748 (n_11391, n12600);
  not g23749 (n_11392, n12615);
  and g23750 (n12616, n_11391, n_11392);
  not g23751 (n_11393, n12616);
  and g23752 (n12617, n_11391, n_11393);
  and g23753 (n12618, n_11392, n_11393);
  not g23754 (n_11394, n12617);
  not g23755 (n_11395, n12618);
  and g23756 (n12619, n_11394, n_11395);
  and g23757 (n12620, n2334, n5666);
  and g23758 (n12621, n2041, n8578);
  and g23759 (n12622, n2331, n6252);
  not g23760 (n_11396, n12621);
  not g23761 (n_11397, n12622);
  and g23762 (n12623, n_11396, n_11397);
  not g23763 (n_11398, n12620);
  not g23764 (n_11399, n12623);
  and g23765 (n12624, n_11398, n_11399);
  not g23766 (n_11400, n12624);
  and g23767 (n12625, \a[48] , n_11400);
  and g23768 (n12626, \a[27] , n12625);
  and g23769 (n12627, n_11398, n_11400);
  and g23770 (n12628, \a[28] , \a[47] );
  and g23771 (n12629, \a[29] , \a[46] );
  not g23772 (n_11401, n12628);
  not g23773 (n_11402, n12629);
  and g23774 (n12630, n_11401, n_11402);
  not g23775 (n_11403, n12630);
  and g23776 (n12631, n12627, n_11403);
  not g23777 (n_11404, n12626);
  not g23778 (n_11405, n12631);
  and g23779 (n12632, n_11404, n_11405);
  not g23780 (n_11406, n12619);
  not g23781 (n_11407, n12632);
  and g23782 (n12633, n_11406, n_11407);
  not g23783 (n_11408, n12633);
  and g23784 (n12634, n_11406, n_11408);
  and g23785 (n12635, n_11407, n_11408);
  not g23786 (n_11409, n12634);
  not g23787 (n_11410, n12635);
  and g23788 (n12636, n_11409, n_11410);
  not g23789 (n_11411, n12636);
  and g23790 (n12637, n12587, n_11411);
  not g23791 (n_11412, n12587);
  and g23792 (n12638, n_11412, n12636);
  and g23793 (n12639, n_11261, n_11264);
  and g23794 (n12640, n12329, n12375);
  not g23795 (n_11413, n12329);
  not g23796 (n_11414, n12375);
  and g23797 (n12641, n_11413, n_11414);
  not g23798 (n_11415, n12640);
  not g23799 (n_11416, n12641);
  and g23800 (n12642, n_11415, n_11416);
  not g23801 (n_11417, n12642);
  and g23802 (n12643, n12281, n_11417);
  not g23803 (n_11418, n12281);
  and g23804 (n12644, n_11418, n12642);
  not g23805 (n_11419, n12643);
  not g23806 (n_11420, n12644);
  and g23807 (n12645, n_11419, n_11420);
  and g23808 (n12646, n_11191, n_11203);
  and g23809 (n12647, n_11154, n_11169);
  and g23810 (n12648, n12646, n12647);
  not g23811 (n_11421, n12646);
  not g23812 (n_11422, n12647);
  and g23813 (n12649, n_11421, n_11422);
  not g23814 (n_11423, n12648);
  not g23815 (n_11424, n12649);
  and g23816 (n12650, n_11423, n_11424);
  and g23817 (n12651, n12645, n12650);
  not g23818 (n_11425, n12645);
  not g23819 (n_11426, n12650);
  and g23820 (n12652, n_11425, n_11426);
  not g23821 (n_11427, n12651);
  not g23822 (n_11428, n12652);
  and g23823 (n12653, n_11427, n_11428);
  not g23824 (n_11429, n12639);
  and g23825 (n12654, n_11429, n12653);
  not g23826 (n_11430, n12653);
  and g23827 (n12655, n12639, n_11430);
  not g23828 (n_11431, n12654);
  not g23829 (n_11432, n12655);
  and g23830 (n12656, n_11431, n_11432);
  not g23831 (n_11433, n12638);
  and g23832 (n12657, n_11433, n12656);
  not g23833 (n_11434, n12637);
  and g23834 (n12658, n_11434, n12657);
  not g23835 (n_11435, n12658);
  and g23836 (n12659, n12656, n_11435);
  and g23837 (n12660, n_11433, n_11435);
  and g23838 (n12661, n_11434, n12660);
  not g23839 (n_11436, n12659);
  not g23840 (n_11437, n12661);
  and g23841 (n12662, n_11436, n_11437);
  not g23842 (n_11438, n12543);
  and g23843 (n12663, n_11438, n12662);
  not g23844 (n_11439, n12662);
  and g23845 (n12664, n12543, n_11439);
  not g23846 (n_11440, n12663);
  not g23847 (n_11441, n12664);
  and g23848 (n12665, n_11440, n_11441);
  and g23849 (n12666, n_11093, n_11097);
  and g23850 (n12667, \a[20] , \a[55] );
  and g23851 (n12668, \a[25] , \a[50] );
  not g23852 (n_11442, n12667);
  not g23853 (n_11443, n12668);
  and g23854 (n12669, n_11442, n_11443);
  and g23855 (n12670, n12667, n12668);
  not g23856 (n_11444, n12670);
  not g23859 (n_11445, n12669);
  not g23861 (n_11446, n12673);
  and g23862 (n12674, n_11444, n_11446);
  and g23863 (n12675, n_11445, n12674);
  and g23864 (n12676, \a[41] , n_11446);
  and g23865 (n12677, \a[34] , n12676);
  not g23866 (n_11447, n12675);
  not g23867 (n_11448, n12677);
  and g23868 (n12678, n_11447, n_11448);
  and g23869 (n12679, n3143, n5018);
  and g23870 (n12680, n2598, n4639);
  and g23871 (n12681, n3812, n5296);
  not g23872 (n_11449, n12680);
  not g23873 (n_11450, n12681);
  and g23874 (n12682, n_11449, n_11450);
  not g23875 (n_11451, n12679);
  not g23876 (n_11452, n12682);
  and g23877 (n12683, n_11451, n_11452);
  not g23878 (n_11453, n12683);
  and g23879 (n12684, \a[44] , n_11453);
  and g23880 (n12685, \a[31] , n12684);
  and g23881 (n12686, \a[33] , \a[42] );
  not g23882 (n_11454, n5294);
  not g23883 (n_11455, n12686);
  and g23884 (n12687, n_11454, n_11455);
  and g23885 (n12688, n_11451, n_11453);
  not g23886 (n_11456, n12687);
  and g23887 (n12689, n_11456, n12688);
  not g23888 (n_11457, n12685);
  not g23889 (n_11458, n12689);
  and g23890 (n12690, n_11457, n_11458);
  not g23891 (n_11459, n12678);
  not g23892 (n_11460, n12690);
  and g23893 (n12691, n_11459, n_11460);
  not g23894 (n_11461, n12691);
  and g23895 (n12692, n_11459, n_11461);
  and g23896 (n12693, n_11460, n_11461);
  not g23897 (n_11462, n12692);
  not g23898 (n_11463, n12693);
  and g23899 (n12694, n_11462, n_11463);
  and g23900 (n12695, n2115, n7232);
  and g23901 (n12696, n1574, n7699);
  and g23902 (n12697, \a[24] , \a[54] );
  and g23903 (n12698, n11867, n12697);
  not g23904 (n_11464, n12696);
  not g23905 (n_11465, n12698);
  and g23906 (n12699, n_11464, n_11465);
  not g23907 (n_11466, n12695);
  not g23908 (n_11467, n12699);
  and g23909 (n12700, n_11466, n_11467);
  not g23910 (n_11468, n12700);
  and g23911 (n12701, \a[54] , n_11468);
  and g23912 (n12702, \a[21] , n12701);
  and g23913 (n12703, n_11466, n_11468);
  and g23914 (n12704, \a[22] , \a[53] );
  and g23915 (n12705, \a[24] , \a[51] );
  not g23916 (n_11469, n12704);
  not g23917 (n_11470, n12705);
  and g23918 (n12706, n_11469, n_11470);
  not g23919 (n_11471, n12706);
  and g23920 (n12707, n12703, n_11471);
  not g23921 (n_11472, n12702);
  not g23922 (n_11473, n12707);
  and g23923 (n12708, n_11472, n_11473);
  not g23924 (n_11474, n12694);
  not g23925 (n_11475, n12708);
  and g23926 (n12709, n_11474, n_11475);
  not g23927 (n_11476, n12709);
  and g23928 (n12710, n_11474, n_11476);
  and g23929 (n12711, n_11475, n_11476);
  not g23930 (n_11477, n12710);
  not g23931 (n_11478, n12711);
  and g23932 (n12712, n_11477, n_11478);
  and g23933 (n12713, n_11233, n_11236);
  not g23934 (n_11479, n12712);
  not g23935 (n_11480, n12713);
  and g23936 (n12714, n_11479, n_11480);
  not g23937 (n_11481, n12714);
  and g23938 (n12715, n_11479, n_11481);
  and g23939 (n12716, n_11480, n_11481);
  not g23940 (n_11482, n12715);
  not g23941 (n_11483, n12716);
  and g23942 (n12717, n_11482, n_11483);
  not g23943 (n_11484, n12666);
  not g23944 (n_11485, n12717);
  and g23945 (n12718, n_11484, n_11485);
  not g23946 (n_11486, n12718);
  and g23947 (n12719, n_11484, n_11486);
  and g23948 (n12720, n_11485, n_11486);
  not g23949 (n_11487, n12719);
  not g23950 (n_11488, n12720);
  and g23951 (n12721, n_11487, n_11488);
  and g23952 (n12722, n_11100, n_11107);
  not g23953 (n_11489, n12721);
  not g23954 (n_11490, n12722);
  and g23955 (n12723, n_11489, n_11490);
  not g23956 (n_11491, n12723);
  and g23957 (n12724, n_11489, n_11491);
  and g23958 (n12725, n_11490, n_11491);
  not g23959 (n_11492, n12724);
  not g23960 (n_11493, n12725);
  and g23961 (n12726, n_11492, n_11493);
  and g23962 (n12727, n_11240, n_11243);
  and g23963 (n12728, n12726, n12727);
  not g23964 (n_11494, n12726);
  not g23965 (n_11495, n12727);
  and g23966 (n12729, n_11494, n_11495);
  not g23967 (n_11496, n12728);
  not g23968 (n_11497, n12729);
  and g23969 (n12730, n_11496, n_11497);
  and g23970 (n12731, n_11246, n_11247);
  not g23971 (n_11498, n12731);
  and g23972 (n12732, n_11108, n_11498);
  not g23973 (n_11499, n12732);
  and g23974 (n12733, n12730, n_11499);
  not g23975 (n_11500, n12730);
  and g23976 (n12734, n_11500, n12732);
  not g23977 (n_11501, n12733);
  not g23978 (n_11502, n12734);
  and g23979 (n12735, n_11501, n_11502);
  and g23980 (n12736, n12665, n12735);
  not g23981 (n_11503, n12665);
  not g23982 (n_11504, n12735);
  and g23983 (n12737, n_11503, n_11504);
  not g23984 (n_11505, n12736);
  not g23985 (n_11506, n12737);
  and g23986 (n12738, n_11505, n_11506);
  not g23987 (n_11507, n12502);
  and g23988 (n12739, n_11507, n12738);
  not g23989 (n_11508, n12738);
  and g23990 (n12740, n12502, n_11508);
  not g23991 (n_11509, n12739);
  not g23992 (n_11510, n12740);
  and g23993 (n12741, n_11509, n_11510);
  and g23994 (n12742, n_11284, n_11288);
  not g23995 (n_11511, n12742);
  and g23996 (n12743, n_11285, n_11511);
  not g23997 (n_11512, n12741);
  and g23998 (n12744, n_11512, n12743);
  not g23999 (n_11513, n12743);
  and g24000 (n12745, n12741, n_11513);
  not g24001 (n_11514, n12744);
  not g24002 (n_11515, n12745);
  and g24003 (\asquared[76] , n_11514, n_11515);
  and g24004 (n12747, n_11510, n_11513);
  not g24005 (n_11516, n12747);
  and g24006 (n12748, n_11509, n_11516);
  and g24007 (n12749, n_11501, n_11505);
  and g24008 (n12750, n_11315, n_11319);
  and g24009 (n12751, n_11416, n_11420);
  and g24010 (n12752, n12750, n12751);
  not g24011 (n_11517, n12750);
  not g24012 (n_11518, n12751);
  and g24013 (n12753, n_11517, n_11518);
  not g24014 (n_11519, n12752);
  not g24015 (n_11520, n12753);
  and g24016 (n12754, n_11519, n_11520);
  and g24017 (n12755, n_11307, n_11311);
  not g24018 (n_11521, n12754);
  and g24019 (n12756, n_11521, n12755);
  not g24020 (n_11522, n12755);
  and g24021 (n12757, n12754, n_11522);
  not g24022 (n_11523, n12756);
  not g24023 (n_11524, n12757);
  and g24024 (n12758, n_11523, n_11524);
  and g24025 (n12759, n_11370, n_11434);
  not g24026 (n_11525, n12759);
  and g24027 (n12760, n12758, n_11525);
  not g24028 (n_11526, n12758);
  and g24029 (n12761, n_11526, n12759);
  not g24030 (n_11527, n12760);
  not g24031 (n_11528, n12761);
  and g24032 (n12762, n_11527, n_11528);
  and g24033 (n12763, n12627, n12674);
  not g24034 (n_11529, n12627);
  not g24035 (n_11530, n12674);
  and g24036 (n12764, n_11529, n_11530);
  not g24037 (n_11531, n12763);
  not g24038 (n_11532, n12764);
  and g24039 (n12765, n_11531, n_11532);
  not g24040 (n_11533, n12765);
  and g24041 (n12766, n12552, n_11533);
  not g24042 (n_11534, n12552);
  and g24043 (n12767, n_11534, n12765);
  not g24044 (n_11535, n12766);
  not g24045 (n_11536, n12767);
  and g24046 (n12768, n_11535, n_11536);
  and g24047 (n12769, n_11461, n_11476);
  and g24048 (n12770, \a[14] , \a[62] );
  not g24049 (n_11537, n12770);
  and g24050 (n12771, n12575, n_11537);
  not g24051 (n_11538, n12575);
  and g24052 (n12772, n_11538, n12770);
  not g24053 (n_11539, n12564);
  not g24054 (n_11540, n12772);
  and g24055 (n12773, n_11539, n_11540);
  not g24056 (n_11541, n12771);
  and g24057 (n12774, n_11541, n12773);
  not g24058 (n_11542, n12774);
  and g24059 (n12775, n_11540, n_11542);
  and g24060 (n12776, n_11541, n12775);
  and g24061 (n12777, n_11539, n_11542);
  not g24062 (n_11543, n12776);
  not g24063 (n_11544, n12777);
  and g24064 (n12778, n_11543, n_11544);
  not g24065 (n_11545, n12769);
  not g24066 (n_11546, n12778);
  and g24067 (n12779, n_11545, n_11546);
  not g24068 (n_11547, n12779);
  and g24069 (n12780, n_11545, n_11547);
  and g24070 (n12781, n_11546, n_11547);
  not g24071 (n_11548, n12780);
  not g24072 (n_11549, n12781);
  and g24073 (n12782, n_11548, n_11549);
  not g24074 (n_11550, n12782);
  and g24075 (n12783, n12768, n_11550);
  not g24076 (n_11551, n12783);
  and g24077 (n12784, n12768, n_11551);
  and g24078 (n12785, n_11550, n_11551);
  not g24079 (n_11552, n12784);
  not g24080 (n_11553, n12785);
  and g24081 (n12786, n_11552, n_11553);
  not g24082 (n_11554, n12786);
  and g24083 (n12787, n12762, n_11554);
  not g24084 (n_11555, n12787);
  and g24085 (n12788, n12762, n_11555);
  and g24086 (n12789, n_11554, n_11555);
  not g24087 (n_11556, n12788);
  not g24088 (n_11557, n12789);
  and g24089 (n12790, n_11556, n_11557);
  and g24090 (n12791, n_11491, n_11497);
  and g24091 (n12792, n12790, n12791);
  not g24092 (n_11558, n12790);
  not g24093 (n_11559, n12791);
  and g24094 (n12793, n_11558, n_11559);
  not g24095 (n_11560, n12792);
  not g24096 (n_11561, n12793);
  and g24097 (n12794, n_11560, n_11561);
  and g24098 (n12795, n_11481, n_11486);
  and g24099 (n12796, n12593, n12610);
  not g24100 (n_11562, n12593);
  not g24101 (n_11563, n12610);
  and g24102 (n12797, n_11562, n_11563);
  not g24103 (n_11564, n12796);
  not g24104 (n_11565, n12797);
  and g24105 (n12798, n_11564, n_11565);
  not g24106 (n_11566, n12798);
  and g24107 (n12799, n12688, n_11566);
  not g24108 (n_11567, n12688);
  and g24109 (n12800, n_11567, n12798);
  not g24110 (n_11568, n12799);
  not g24111 (n_11569, n12800);
  and g24112 (n12801, n_11568, n_11569);
  and g24113 (n12802, n_11393, n_11408);
  and g24114 (n12803, n_11352, n_11364);
  and g24115 (n12804, n12802, n12803);
  not g24116 (n_11570, n12802);
  not g24117 (n_11571, n12803);
  and g24118 (n12805, n_11570, n_11571);
  not g24119 (n_11572, n12804);
  not g24120 (n_11573, n12805);
  and g24121 (n12806, n_11572, n_11573);
  and g24122 (n12807, n12801, n12806);
  not g24123 (n_11574, n12801);
  not g24124 (n_11575, n12806);
  and g24125 (n12808, n_11574, n_11575);
  not g24126 (n_11576, n12807);
  not g24127 (n_11577, n12808);
  and g24128 (n12809, n_11576, n_11577);
  not g24129 (n_11578, n12809);
  and g24130 (n12810, n12795, n_11578);
  not g24131 (n_11579, n12795);
  and g24132 (n12811, n_11579, n12809);
  not g24133 (n_11580, n12810);
  not g24134 (n_11581, n12811);
  and g24135 (n12812, n_11580, n_11581);
  and g24136 (n12813, n2617, n5666);
  and g24137 (n12814, n3110, n8578);
  and g24138 (n12815, n2334, n6252);
  not g24139 (n_11582, n12814);
  not g24140 (n_11583, n12815);
  and g24141 (n12816, n_11582, n_11583);
  not g24142 (n_11584, n12813);
  not g24143 (n_11585, n12816);
  and g24144 (n12817, n_11584, n_11585);
  not g24145 (n_11586, n12817);
  and g24146 (n12818, n_11584, n_11586);
  and g24147 (n12819, \a[29] , \a[47] );
  and g24148 (n12820, \a[30] , \a[46] );
  not g24149 (n_11587, n12819);
  not g24150 (n_11588, n12820);
  and g24151 (n12821, n_11587, n_11588);
  not g24152 (n_11589, n12821);
  and g24153 (n12822, n12818, n_11589);
  and g24154 (n12823, \a[48] , n_11586);
  and g24155 (n12824, \a[28] , n12823);
  not g24156 (n_11590, n12822);
  not g24157 (n_11591, n12824);
  and g24158 (n12825, n_11590, n_11591);
  and g24159 (n12826, n3828, n5413);
  and g24160 (n12827, n4595, n6453);
  and g24161 (n12828, n3319, n5344);
  not g24162 (n_11592, n12827);
  not g24163 (n_11593, n12828);
  and g24164 (n12829, n_11592, n_11593);
  not g24165 (n_11594, n12826);
  not g24166 (n_11595, n12829);
  and g24167 (n12830, n_11594, n_11595);
  not g24168 (n_11596, n12830);
  and g24169 (n12831, \a[42] , n_11596);
  and g24170 (n12832, \a[34] , n12831);
  and g24171 (n12833, n_11594, n_11596);
  and g24172 (n12834, \a[35] , \a[41] );
  and g24173 (n12835, \a[36] , \a[40] );
  not g24174 (n_11597, n12834);
  not g24175 (n_11598, n12835);
  and g24176 (n12836, n_11597, n_11598);
  not g24177 (n_11599, n12836);
  and g24178 (n12837, n12833, n_11599);
  not g24179 (n_11600, n12832);
  not g24180 (n_11601, n12837);
  and g24181 (n12838, n_11600, n_11601);
  not g24182 (n_11602, n12825);
  not g24183 (n_11603, n12838);
  and g24184 (n12839, n_11602, n_11603);
  not g24185 (n_11604, n12839);
  and g24186 (n12840, n_11602, n_11604);
  and g24187 (n12841, n_11603, n_11604);
  not g24188 (n_11605, n12840);
  not g24189 (n_11606, n12841);
  and g24190 (n12842, n_11605, n_11606);
  and g24191 (n12843, \a[24] , \a[52] );
  and g24192 (n12844, \a[25] , \a[51] );
  not g24193 (n_11607, n12843);
  not g24194 (n_11608, n12844);
  and g24195 (n12845, n_11607, n_11608);
  and g24196 (n12846, n1904, n6968);
  not g24197 (n_11609, n12846);
  and g24198 (n12847, n5430, n_11609);
  not g24199 (n_11610, n12845);
  and g24200 (n12848, n_11610, n12847);
  not g24201 (n_11611, n12848);
  and g24202 (n12849, n5430, n_11611);
  and g24203 (n12850, n_11609, n_11611);
  and g24204 (n12851, n_11610, n12850);
  not g24205 (n_11612, n12849);
  not g24206 (n_11613, n12851);
  and g24207 (n12852, n_11612, n_11613);
  not g24208 (n_11614, n12842);
  not g24209 (n_11615, n12852);
  and g24210 (n12853, n_11614, n_11615);
  not g24211 (n_11616, n12853);
  and g24212 (n12854, n_11614, n_11616);
  and g24213 (n12855, n_11615, n_11616);
  not g24214 (n_11617, n12854);
  not g24215 (n_11618, n12855);
  and g24216 (n12856, n_11617, n_11618);
  and g24217 (n12857, n_11294, n_11298);
  and g24218 (n12858, n12856, n12857);
  not g24219 (n_11619, n12856);
  not g24220 (n_11620, n12857);
  and g24221 (n12859, n_11619, n_11620);
  not g24222 (n_11621, n12858);
  not g24223 (n_11622, n12859);
  and g24224 (n12860, n_11621, n_11622);
  and g24225 (n12861, n1048, n9509);
  and g24226 (n12862, n993, n8905);
  and g24227 (n12863, n891, n9512);
  not g24228 (n_11623, n12862);
  not g24229 (n_11624, n12863);
  and g24230 (n12864, n_11623, n_11624);
  not g24231 (n_11625, n12861);
  not g24232 (n_11626, n12864);
  and g24233 (n12865, n_11625, n_11626);
  not g24234 (n_11627, n12865);
  and g24235 (n12866, \a[61] , n_11627);
  and g24236 (n12867, \a[15] , n12866);
  and g24237 (n12868, n_11625, n_11627);
  and g24238 (n12869, \a[16] , \a[60] );
  and g24239 (n12870, \a[17] , \a[59] );
  not g24240 (n_11628, n12869);
  not g24241 (n_11629, n12870);
  and g24242 (n12871, n_11628, n_11629);
  not g24243 (n_11630, n12871);
  and g24244 (n12872, n12868, n_11630);
  not g24245 (n_11631, n12867);
  not g24246 (n_11632, n12872);
  and g24247 (n12873, n_11631, n_11632);
  not g24248 (n_11633, n12873);
  and g24249 (n12874, n12703, n_11633);
  not g24250 (n_11634, n12703);
  and g24251 (n12875, n_11634, n12873);
  not g24252 (n_11635, n12874);
  not g24253 (n_11636, n12875);
  and g24254 (n12876, n_11635, n_11636);
  and g24255 (n12877, \a[26] , \a[50] );
  and g24256 (n12878, \a[27] , \a[49] );
  not g24257 (n_11637, n12877);
  not g24258 (n_11638, n12878);
  and g24259 (n12879, n_11637, n_11638);
  and g24260 (n12880, n2227, n6325);
  not g24261 (n_11639, n12880);
  not g24264 (n_11640, n12879);
  not g24266 (n_11641, n12883);
  and g24267 (n12884, \a[58] , n_11641);
  and g24268 (n12885, \a[18] , n12884);
  and g24269 (n12886, n_11639, n_11641);
  and g24270 (n12887, n_11640, n12886);
  not g24271 (n_11642, n12885);
  not g24272 (n_11643, n12887);
  and g24273 (n12888, n_11642, n_11643);
  not g24274 (n_11644, n12876);
  not g24275 (n_11645, n12888);
  and g24276 (n12889, n_11644, n_11645);
  and g24277 (n12890, n12876, n12888);
  not g24278 (n_11646, n12889);
  not g24279 (n_11647, n12890);
  and g24280 (n12891, n_11646, n_11647);
  and g24281 (n12892, n12860, n12891);
  not g24282 (n_11648, n12860);
  not g24283 (n_11649, n12891);
  and g24284 (n12893, n_11648, n_11649);
  not g24285 (n_11650, n12893);
  and g24286 (n12894, n12812, n_11650);
  not g24287 (n_11651, n12892);
  and g24288 (n12895, n_11651, n12894);
  not g24289 (n_11652, n12895);
  and g24290 (n12896, n12812, n_11652);
  and g24291 (n12897, n_11650, n_11652);
  and g24292 (n12898, n_11651, n12897);
  not g24293 (n_11653, n12896);
  not g24294 (n_11654, n12898);
  and g24295 (n12899, n_11653, n_11654);
  not g24296 (n_11655, n12899);
  and g24297 (n12900, n12794, n_11655);
  not g24298 (n_11656, n12794);
  and g24299 (n12901, n_11656, n12899);
  and g24300 (n12902, n_11335, n_11441);
  and g24301 (n12903, n_11431, n_11435);
  and g24302 (n12904, n_11302, n_11330);
  and g24303 (n12905, n_11322, n_11326);
  and g24304 (n12906, \a[31] , \a[45] );
  and g24305 (n12907, \a[32] , \a[44] );
  not g24306 (n_11657, n12906);
  not g24307 (n_11658, n12907);
  and g24308 (n12908, n_11657, n_11658);
  and g24309 (n12909, n3812, n5713);
  not g24310 (n_11659, n12909);
  not g24312 (n_11660, n12908);
  not g24315 (n_11661, n12912);
  and g24316 (n12913, n_11659, n_11661);
  and g24317 (n12914, n_11660, n12913);
  and g24318 (n12915, \a[63] , n_11661);
  and g24319 (n12916, \a[13] , n12915);
  not g24320 (n_11662, n12914);
  not g24321 (n_11663, n12916);
  and g24322 (n12917, n_11662, n_11663);
  and g24323 (n12918, \a[19] , \a[57] );
  and g24324 (n12919, \a[23] , \a[53] );
  not g24325 (n_11664, n12918);
  not g24326 (n_11665, n12919);
  and g24327 (n12920, n_11664, n_11665);
  and g24328 (n12921, n12918, n12919);
  not g24329 (n_11666, n12921);
  and g24330 (n12922, n5449, n_11666);
  not g24331 (n_11667, n12920);
  and g24332 (n12923, n_11667, n12922);
  not g24333 (n_11668, n12923);
  and g24334 (n12924, n5449, n_11668);
  and g24335 (n12925, n_11666, n_11668);
  and g24336 (n12926, n_11667, n12925);
  not g24337 (n_11669, n12924);
  not g24338 (n_11670, n12926);
  and g24339 (n12927, n_11669, n_11670);
  not g24340 (n_11671, n12917);
  not g24341 (n_11672, n12927);
  and g24342 (n12928, n_11671, n_11672);
  not g24343 (n_11673, n12928);
  and g24344 (n12929, n_11671, n_11673);
  and g24345 (n12930, n_11672, n_11673);
  not g24346 (n_11674, n12929);
  not g24347 (n_11675, n12930);
  and g24348 (n12931, n_11674, n_11675);
  and g24349 (n12932, n1574, n7701);
  and g24350 (n12933, n1693, n7421);
  and g24351 (n12934, n1494, n9161);
  not g24352 (n_11676, n12933);
  not g24353 (n_11677, n12934);
  and g24354 (n12935, n_11676, n_11677);
  not g24355 (n_11678, n12932);
  not g24356 (n_11679, n12935);
  and g24357 (n12936, n_11678, n_11679);
  not g24358 (n_11680, n12936);
  and g24359 (n12937, n9985, n_11680);
  and g24360 (n12938, n_11678, n_11680);
  and g24361 (n12939, \a[21] , \a[55] );
  and g24362 (n12940, \a[22] , \a[54] );
  not g24363 (n_11681, n12939);
  not g24364 (n_11682, n12940);
  and g24365 (n12941, n_11681, n_11682);
  not g24366 (n_11683, n12941);
  and g24367 (n12942, n12938, n_11683);
  not g24368 (n_11684, n12937);
  not g24369 (n_11685, n12942);
  and g24370 (n12943, n_11684, n_11685);
  not g24371 (n_11686, n12931);
  not g24372 (n_11687, n12943);
  and g24373 (n12944, n_11686, n_11687);
  not g24374 (n_11688, n12944);
  and g24375 (n12945, n_11686, n_11688);
  and g24376 (n12946, n_11687, n_11688);
  not g24377 (n_11689, n12945);
  not g24378 (n_11690, n12946);
  and g24379 (n12947, n_11689, n_11690);
  and g24380 (n12948, n_11424, n_11427);
  not g24381 (n_11691, n12947);
  not g24382 (n_11692, n12948);
  and g24383 (n12949, n_11691, n_11692);
  and g24384 (n12950, n12947, n12948);
  not g24385 (n_11693, n12949);
  not g24386 (n_11694, n12950);
  and g24387 (n12951, n_11693, n_11694);
  not g24388 (n_11695, n12905);
  and g24389 (n12952, n_11695, n12951);
  not g24390 (n_11696, n12951);
  and g24391 (n12953, n12905, n_11696);
  not g24392 (n_11697, n12952);
  not g24393 (n_11698, n12953);
  and g24394 (n12954, n_11697, n_11698);
  not g24395 (n_11699, n12904);
  and g24396 (n12955, n_11699, n12954);
  not g24397 (n_11700, n12954);
  and g24398 (n12956, n12904, n_11700);
  not g24399 (n_11701, n12955);
  not g24400 (n_11702, n12956);
  and g24401 (n12957, n_11701, n_11702);
  not g24402 (n_11703, n12903);
  and g24403 (n12958, n_11703, n12957);
  not g24404 (n_11704, n12957);
  and g24405 (n12959, n12903, n_11704);
  not g24406 (n_11705, n12958);
  not g24407 (n_11706, n12959);
  and g24408 (n12960, n_11705, n_11706);
  not g24409 (n_11707, n12902);
  and g24410 (n12961, n_11707, n12960);
  not g24411 (n_11708, n12960);
  and g24412 (n12962, n12902, n_11708);
  not g24413 (n_11709, n12961);
  not g24414 (n_11710, n12962);
  and g24415 (n12963, n_11709, n_11710);
  not g24416 (n_11711, n12901);
  and g24417 (n12964, n_11711, n12963);
  not g24418 (n_11712, n12900);
  and g24419 (n12965, n_11712, n12964);
  not g24420 (n_11713, n12965);
  and g24421 (n12966, n12963, n_11713);
  and g24422 (n12967, n_11711, n_11713);
  and g24423 (n12968, n_11712, n12967);
  not g24424 (n_11714, n12966);
  not g24425 (n_11715, n12968);
  and g24426 (n12969, n_11714, n_11715);
  not g24427 (n_11716, n12749);
  not g24428 (n_11717, n12969);
  and g24429 (n12970, n_11716, n_11717);
  and g24430 (n12971, n12749, n12969);
  not g24431 (n_11718, n12970);
  not g24432 (n_11719, n12971);
  and g24433 (n12972, n_11718, n_11719);
  not g24434 (n_11720, n12748);
  and g24435 (n12973, n_11720, n12972);
  not g24436 (n_11721, n12972);
  and g24437 (n12974, n12748, n_11721);
  not g24438 (n_11722, n12973);
  not g24439 (n_11723, n12974);
  and g24440 (\asquared[77] , n_11722, n_11723);
  and g24441 (n12976, n_11709, n_11713);
  and g24442 (n12977, n_11701, n_11705);
  and g24443 (n12978, n1052, n9509);
  not g24444 (n_11724, n12978);
  and g24445 (n12979, \a[59] , n_11724);
  and g24446 (n12980, \a[18] , n12979);
  and g24447 (n12981, \a[60] , n_11724);
  and g24448 (n12982, \a[17] , n12981);
  not g24449 (n_11725, n12980);
  not g24450 (n_11726, n12982);
  and g24451 (n12983, n_11725, n_11726);
  not g24452 (n_11727, n12850);
  not g24453 (n_11728, n12983);
  and g24454 (n12984, n_11727, n_11728);
  not g24455 (n_11729, n12984);
  and g24456 (n12985, n_11727, n_11729);
  and g24457 (n12986, n_11728, n_11729);
  not g24458 (n_11730, n12985);
  not g24459 (n_11731, n12986);
  and g24460 (n12987, n_11730, n_11731);
  and g24461 (n12988, n_11565, n_11569);
  and g24462 (n12989, n12987, n12988);
  not g24463 (n_11732, n12987);
  not g24464 (n_11733, n12988);
  and g24465 (n12990, n_11732, n_11733);
  not g24466 (n_11734, n12989);
  not g24467 (n_11735, n12990);
  and g24468 (n12991, n_11734, n_11735);
  and g24469 (n12992, n_11532, n_11536);
  not g24470 (n_11736, n12991);
  and g24471 (n12993, n_11736, n12992);
  not g24472 (n_11737, n12992);
  and g24473 (n12994, n12991, n_11737);
  not g24474 (n_11738, n12993);
  not g24475 (n_11739, n12994);
  and g24476 (n12995, n_11738, n_11739);
  and g24477 (n12996, n_11622, n_11651);
  not g24478 (n_11740, n12996);
  and g24479 (n12997, n12995, n_11740);
  not g24480 (n_11741, n12995);
  and g24481 (n12998, n_11741, n12996);
  not g24482 (n_11742, n12997);
  not g24483 (n_11743, n12998);
  and g24484 (n12999, n_11742, n_11743);
  and g24485 (n13000, n12818, n12938);
  not g24486 (n_11744, n12818);
  not g24487 (n_11745, n12938);
  and g24488 (n13001, n_11744, n_11745);
  not g24489 (n_11746, n13000);
  not g24490 (n_11747, n13001);
  and g24491 (n13002, n_11746, n_11747);
  not g24492 (n_11748, n13002);
  and g24493 (n13003, n12913, n_11748);
  not g24494 (n_11749, n12913);
  and g24495 (n13004, n_11749, n13002);
  not g24496 (n_11750, n13003);
  not g24497 (n_11751, n13004);
  and g24498 (n13005, n_11750, n_11751);
  and g24499 (n13006, n12868, n12886);
  not g24500 (n_11752, n12868);
  not g24501 (n_11753, n12886);
  and g24502 (n13007, n_11752, n_11753);
  not g24503 (n_11754, n13006);
  not g24504 (n_11755, n13007);
  and g24505 (n13008, n_11754, n_11755);
  not g24506 (n_11756, n13008);
  and g24507 (n13009, n12925, n_11756);
  not g24508 (n_11757, n12925);
  and g24509 (n13010, n_11757, n13008);
  not g24510 (n_11758, n13009);
  not g24511 (n_11759, n13010);
  and g24512 (n13011, n_11758, n_11759);
  and g24513 (n13012, n_11673, n_11688);
  not g24514 (n_11760, n13011);
  and g24515 (n13013, n_11760, n13012);
  not g24516 (n_11761, n13012);
  and g24517 (n13014, n13011, n_11761);
  not g24518 (n_11762, n13013);
  not g24519 (n_11763, n13014);
  and g24520 (n13015, n_11762, n_11763);
  and g24521 (n13016, n13005, n13015);
  not g24522 (n_11764, n13005);
  not g24523 (n_11765, n13015);
  and g24524 (n13017, n_11764, n_11765);
  not g24525 (n_11766, n13016);
  not g24526 (n_11767, n13017);
  and g24527 (n13018, n_11766, n_11767);
  and g24528 (n13019, n12999, n13018);
  not g24529 (n_11768, n12999);
  not g24530 (n_11769, n13018);
  and g24531 (n13020, n_11768, n_11769);
  not g24532 (n_11770, n13019);
  not g24533 (n_11771, n13020);
  and g24534 (n13021, n_11770, n_11771);
  not g24535 (n_11772, n13021);
  and g24536 (n13022, n12977, n_11772);
  not g24537 (n_11773, n12977);
  and g24538 (n13023, n_11773, n13021);
  not g24539 (n_11774, n13022);
  not g24540 (n_11775, n13023);
  and g24541 (n13024, n_11774, n_11775);
  and g24542 (n13025, n_11634, n_11633);
  not g24543 (n_11776, n13025);
  and g24544 (n13026, n_11646, n_11776);
  and g24545 (n13027, n12775, n13026);
  not g24546 (n_11777, n12775);
  not g24547 (n_11778, n13026);
  and g24548 (n13028, n_11777, n_11778);
  not g24549 (n_11779, n13027);
  not g24550 (n_11780, n13028);
  and g24551 (n13029, n_11779, n_11780);
  and g24552 (n13030, n_11604, n_11616);
  not g24553 (n_11781, n13029);
  and g24554 (n13031, n_11781, n13030);
  not g24555 (n_11782, n13030);
  and g24556 (n13032, n13029, n_11782);
  not g24557 (n_11783, n13031);
  not g24558 (n_11784, n13032);
  and g24559 (n13033, n_11783, n_11784);
  and g24560 (n13034, n_11693, n_11697);
  not g24561 (n_11785, n13033);
  and g24562 (n13035, n_11785, n13034);
  not g24563 (n_11786, n13034);
  and g24564 (n13036, n13033, n_11786);
  not g24565 (n_11787, n13035);
  not g24566 (n_11788, n13036);
  and g24567 (n13037, n_11787, n_11788);
  and g24568 (n13038, \a[31] , \a[63] );
  and g24569 (n13039, n7400, n13038);
  and g24570 (n13040, n2865, n5666);
  and g24571 (n13041, \a[14] , \a[63] );
  and g24572 (n13042, \a[30] , \a[47] );
  and g24573 (n13043, n13041, n13042);
  not g24574 (n_11789, n13040);
  not g24575 (n_11790, n13043);
  and g24576 (n13044, n_11789, n_11790);
  not g24577 (n_11791, n13039);
  not g24578 (n_11792, n13044);
  and g24579 (n13045, n_11791, n_11792);
  not g24580 (n_11793, n13045);
  and g24581 (n13046, n_11791, n_11793);
  and g24582 (n13047, \a[31] , \a[46] );
  not g24583 (n_11794, n13041);
  not g24584 (n_11795, n13047);
  and g24585 (n13048, n_11794, n_11795);
  not g24586 (n_11796, n13048);
  and g24587 (n13049, n13046, n_11796);
  and g24588 (n13050, n13042, n_11793);
  not g24589 (n_11797, n13049);
  not g24590 (n_11798, n13050);
  and g24591 (n13051, n_11797, n_11798);
  and g24592 (n13052, \a[35] , \a[42] );
  and g24593 (n13053, n3687, n5413);
  and g24594 (n13054, n5031, n6453);
  and g24595 (n13055, n3828, n5344);
  not g24596 (n_11799, n13054);
  not g24597 (n_11800, n13055);
  and g24598 (n13056, n_11799, n_11800);
  not g24599 (n_11801, n13053);
  not g24600 (n_11802, n13056);
  and g24601 (n13057, n_11801, n_11802);
  not g24602 (n_11803, n13057);
  and g24603 (n13058, n13052, n_11803);
  and g24604 (n13059, n_11801, n_11803);
  and g24605 (n13060, \a[36] , \a[41] );
  not g24606 (n_11804, n5695);
  not g24607 (n_11805, n13060);
  and g24608 (n13061, n_11804, n_11805);
  not g24609 (n_11806, n13061);
  and g24610 (n13062, n13059, n_11806);
  not g24611 (n_11807, n13058);
  not g24612 (n_11808, n13062);
  and g24613 (n13063, n_11807, n_11808);
  not g24614 (n_11809, n13051);
  not g24615 (n_11810, n13063);
  and g24616 (n13064, n_11809, n_11810);
  not g24617 (n_11811, n13064);
  and g24618 (n13065, n_11809, n_11811);
  and g24619 (n13066, n_11810, n_11811);
  not g24620 (n_11812, n13065);
  not g24621 (n_11813, n13066);
  and g24622 (n13067, n_11812, n_11813);
  and g24623 (n13068, \a[62] , n6981);
  not g24624 (n_11814, n13068);
  and g24625 (n13069, n5083, n_11814);
  not g24626 (n_11815, n13069);
  and g24627 (n13070, n5083, n_11815);
  and g24628 (n13071, n_11814, n_11815);
  and g24629 (n13072, \a[15] , \a[62] );
  not g24630 (n_11816, \a[39] );
  not g24631 (n_11817, n13072);
  and g24632 (n13073, n_11816, n_11817);
  not g24633 (n_11818, n13073);
  and g24634 (n13074, n13071, n_11818);
  not g24635 (n_11819, n13070);
  not g24636 (n_11820, n13074);
  and g24637 (n13075, n_11819, n_11820);
  not g24638 (n_11821, n13067);
  not g24639 (n_11822, n13075);
  and g24640 (n13076, n_11821, n_11822);
  not g24641 (n_11823, n13076);
  and g24642 (n13077, n_11821, n_11823);
  and g24643 (n13078, n_11822, n_11823);
  not g24644 (n_11824, n13077);
  not g24645 (n_11825, n13078);
  and g24646 (n13079, n_11824, n_11825);
  and g24647 (n13080, n_11520, n_11524);
  and g24648 (n13081, n13079, n13080);
  not g24649 (n_11826, n13079);
  not g24650 (n_11827, n13080);
  and g24651 (n13082, n_11826, n_11827);
  not g24652 (n_11828, n13081);
  not g24653 (n_11829, n13082);
  and g24654 (n13083, n_11828, n_11829);
  and g24655 (n13084, n1494, n8200);
  and g24656 (n13085, n1492, n7942);
  and g24657 (n13086, n1490, n8436);
  not g24658 (n_11830, n13085);
  not g24659 (n_11831, n13086);
  and g24660 (n13087, n_11830, n_11831);
  not g24661 (n_11832, n13084);
  not g24662 (n_11833, n13087);
  and g24663 (n13088, n_11832, n_11833);
  not g24664 (n_11834, n13088);
  and g24665 (n13089, \a[58] , n_11834);
  and g24666 (n13090, \a[19] , n13089);
  and g24667 (n13091, n_11832, n_11834);
  and g24668 (n13092, \a[21] , \a[56] );
  not g24669 (n_11835, n10658);
  not g24670 (n_11836, n13092);
  and g24671 (n13093, n_11835, n_11836);
  not g24672 (n_11837, n13093);
  and g24673 (n13094, n13091, n_11837);
  not g24674 (n_11838, n13090);
  not g24675 (n_11839, n13094);
  and g24676 (n13095, n_11838, n_11839);
  not g24677 (n_11840, n13095);
  and g24678 (n13096, n12833, n_11840);
  not g24679 (n_11841, n12833);
  and g24680 (n13097, n_11841, n13095);
  not g24681 (n_11842, n13096);
  not g24682 (n_11843, n13097);
  and g24683 (n13098, n_11842, n_11843);
  and g24684 (n13099, n2334, n6256);
  and g24685 (n13100, n2041, n5888);
  and g24686 (n13101, n2331, n6325);
  not g24687 (n_11844, n13100);
  not g24688 (n_11845, n13101);
  and g24689 (n13102, n_11844, n_11845);
  not g24690 (n_11846, n13099);
  not g24691 (n_11847, n13102);
  and g24692 (n13103, n_11846, n_11847);
  not g24693 (n_11848, n13103);
  and g24694 (n13104, \a[50] , n_11848);
  and g24695 (n13105, \a[27] , n13104);
  and g24696 (n13106, n_11846, n_11848);
  and g24697 (n13107, \a[28] , \a[49] );
  and g24698 (n13108, \a[29] , \a[48] );
  not g24699 (n_11849, n13107);
  not g24700 (n_11850, n13108);
  and g24701 (n13109, n_11849, n_11850);
  not g24702 (n_11851, n13109);
  and g24703 (n13110, n13106, n_11851);
  not g24704 (n_11852, n13105);
  not g24705 (n_11853, n13110);
  and g24706 (n13111, n_11852, n_11853);
  not g24707 (n_11854, n13098);
  not g24708 (n_11855, n13111);
  and g24709 (n13112, n_11854, n_11855);
  and g24710 (n13113, n13098, n13111);
  not g24711 (n_11856, n13112);
  not g24712 (n_11857, n13113);
  and g24713 (n13114, n_11856, n_11857);
  and g24714 (n13115, n13083, n13114);
  not g24715 (n_11858, n13083);
  not g24716 (n_11859, n13114);
  and g24717 (n13116, n_11858, n_11859);
  not g24718 (n_11860, n13116);
  and g24719 (n13117, n13037, n_11860);
  not g24720 (n_11861, n13115);
  and g24721 (n13118, n_11861, n13117);
  not g24722 (n_11862, n13118);
  and g24723 (n13119, n13037, n_11862);
  and g24724 (n13120, n_11860, n_11862);
  and g24725 (n13121, n_11861, n13120);
  not g24726 (n_11863, n13119);
  not g24727 (n_11864, n13121);
  and g24728 (n13122, n_11863, n_11864);
  not g24729 (n_11865, n13122);
  and g24730 (n13123, n13024, n_11865);
  not g24731 (n_11866, n13024);
  and g24732 (n13124, n_11866, n13122);
  and g24733 (n13125, n_11561, n_11712);
  and g24734 (n13126, n_11581, n_11652);
  and g24735 (n13127, n_11527, n_11555);
  and g24736 (n13128, n_11547, n_11551);
  and g24737 (n13129, \a[22] , \a[55] );
  and g24738 (n13130, \a[26] , \a[51] );
  not g24739 (n_11867, n13129);
  not g24740 (n_11868, n13130);
  and g24741 (n13131, n_11867, n_11868);
  and g24742 (n13132, n13129, n13130);
  not g24743 (n_11869, n13132);
  not g24746 (n_11870, n13131);
  not g24748 (n_11871, n13135);
  and g24749 (n13136, n_11869, n_11871);
  and g24750 (n13137, n_11870, n13136);
  and g24751 (n13138, \a[43] , n_11871);
  and g24752 (n13139, \a[34] , n13138);
  not g24753 (n_11872, n13137);
  not g24754 (n_11873, n13139);
  and g24755 (n13140, n_11872, n_11873);
  and g24756 (n13141, n1666, n7699);
  and g24757 (n13142, n1547, n10905);
  and g24758 (n13143, n1904, n7433);
  not g24759 (n_11874, n13142);
  not g24760 (n_11875, n13143);
  and g24761 (n13144, n_11874, n_11875);
  not g24762 (n_11876, n13141);
  not g24763 (n_11877, n13144);
  and g24764 (n13145, n_11876, n_11877);
  not g24765 (n_11878, n13145);
  and g24766 (n13146, \a[52] , n_11878);
  and g24767 (n13147, \a[25] , n13146);
  and g24768 (n13148, \a[23] , \a[54] );
  and g24769 (n13149, \a[24] , \a[53] );
  not g24770 (n_11879, n13148);
  not g24771 (n_11880, n13149);
  and g24772 (n13150, n_11879, n_11880);
  and g24773 (n13151, n_11876, n_11878);
  not g24774 (n_11881, n13150);
  and g24775 (n13152, n_11881, n13151);
  not g24776 (n_11882, n13147);
  not g24777 (n_11883, n13152);
  and g24778 (n13153, n_11882, n_11883);
  not g24779 (n_11884, n13140);
  not g24780 (n_11885, n13153);
  and g24781 (n13154, n_11884, n_11885);
  not g24782 (n_11886, n13154);
  and g24783 (n13155, n_11884, n_11886);
  and g24784 (n13156, n_11885, n_11886);
  not g24785 (n_11887, n13155);
  not g24786 (n_11888, n13156);
  and g24787 (n13157, n_11887, n_11888);
  and g24788 (n13158, \a[32] , \a[45] );
  not g24789 (n_11889, n5451);
  not g24790 (n_11890, n13158);
  and g24791 (n13159, n_11889, n_11890);
  and g24792 (n13160, n3143, n5713);
  not g24793 (n_11891, n13160);
  not g24796 (n_11892, n13159);
  not g24798 (n_11893, n13163);
  and g24799 (n13164, \a[61] , n_11893);
  and g24800 (n13165, \a[16] , n13164);
  and g24801 (n13166, n_11891, n_11893);
  and g24802 (n13167, n_11892, n13166);
  not g24803 (n_11894, n13165);
  not g24804 (n_11895, n13167);
  and g24805 (n13168, n_11894, n_11895);
  not g24806 (n_11896, n13157);
  not g24807 (n_11897, n13168);
  and g24808 (n13169, n_11896, n_11897);
  not g24809 (n_11898, n13169);
  and g24810 (n13170, n_11896, n_11898);
  and g24811 (n13171, n_11897, n_11898);
  not g24812 (n_11899, n13170);
  not g24813 (n_11900, n13171);
  and g24814 (n13172, n_11899, n_11900);
  and g24815 (n13173, n_11573, n_11576);
  not g24816 (n_11901, n13172);
  not g24817 (n_11902, n13173);
  and g24818 (n13174, n_11901, n_11902);
  not g24819 (n_11903, n13174);
  and g24820 (n13175, n_11901, n_11903);
  and g24821 (n13176, n_11902, n_11903);
  not g24822 (n_11904, n13175);
  not g24823 (n_11905, n13176);
  and g24824 (n13177, n_11904, n_11905);
  not g24825 (n_11906, n13128);
  not g24826 (n_11907, n13177);
  and g24827 (n13178, n_11906, n_11907);
  and g24828 (n13179, n13128, n_11905);
  and g24829 (n13180, n_11904, n13179);
  not g24830 (n_11908, n13178);
  not g24831 (n_11909, n13180);
  and g24832 (n13181, n_11908, n_11909);
  not g24833 (n_11910, n13127);
  and g24834 (n13182, n_11910, n13181);
  not g24835 (n_11911, n13181);
  and g24836 (n13183, n13127, n_11911);
  not g24837 (n_11912, n13182);
  not g24838 (n_11913, n13183);
  and g24839 (n13184, n_11912, n_11913);
  not g24840 (n_11914, n13126);
  and g24841 (n13185, n_11914, n13184);
  not g24842 (n_11915, n13184);
  and g24843 (n13186, n13126, n_11915);
  not g24844 (n_11916, n13185);
  not g24845 (n_11917, n13186);
  and g24846 (n13187, n_11916, n_11917);
  not g24847 (n_11918, n13125);
  and g24848 (n13188, n_11918, n13187);
  not g24849 (n_11919, n13187);
  and g24850 (n13189, n13125, n_11919);
  not g24851 (n_11920, n13188);
  not g24852 (n_11921, n13189);
  and g24853 (n13190, n_11920, n_11921);
  not g24854 (n_11922, n13124);
  and g24855 (n13191, n_11922, n13190);
  not g24856 (n_11923, n13123);
  and g24857 (n13192, n_11923, n13191);
  not g24858 (n_11924, n13192);
  and g24859 (n13193, n13190, n_11924);
  and g24860 (n13194, n_11922, n_11924);
  and g24861 (n13195, n_11923, n13194);
  not g24862 (n_11925, n13193);
  not g24863 (n_11926, n13195);
  and g24864 (n13196, n_11925, n_11926);
  not g24865 (n_11927, n12976);
  not g24866 (n_11928, n13196);
  and g24867 (n13197, n_11927, n_11928);
  and g24868 (n13198, n12976, n13196);
  not g24869 (n_11929, n13197);
  not g24870 (n_11930, n13198);
  and g24871 (n13199, n_11929, n_11930);
  and g24872 (n13200, n_11720, n_11719);
  not g24873 (n_11931, n13200);
  and g24874 (n13201, n_11718, n_11931);
  not g24875 (n_11932, n13199);
  and g24876 (n13202, n_11932, n13201);
  not g24877 (n_11933, n13201);
  and g24878 (n13203, n13199, n_11933);
  not g24879 (n_11934, n13202);
  not g24880 (n_11935, n13203);
  and g24881 (\asquared[78] , n_11934, n_11935);
  and g24882 (n13205, n_11930, n_11933);
  not g24883 (n_11936, n13205);
  and g24884 (n13206, n_11929, n_11936);
  and g24885 (n13207, n_11920, n_11924);
  and g24886 (n13208, n_11788, n_11862);
  and g24887 (n13209, n_11742, n_11770);
  and g24888 (n13210, n_11780, n_11784);
  and g24889 (n13211, n1492, n8985);
  and g24890 (n13212, \a[57] , \a[60] );
  and g24891 (n13213, n3648, n13212);
  and g24892 (n13214, n1149, n9509);
  not g24893 (n_11937, n13213);
  not g24894 (n_11938, n13214);
  and g24895 (n13215, n_11937, n_11938);
  not g24896 (n_11939, n13211);
  not g24897 (n_11940, n13215);
  and g24898 (n13216, n_11939, n_11940);
  not g24899 (n_11941, n13216);
  and g24900 (n13217, n_11939, n_11941);
  and g24901 (n13218, \a[19] , \a[59] );
  and g24902 (n13219, \a[21] , \a[57] );
  not g24903 (n_11942, n13218);
  not g24904 (n_11943, n13219);
  and g24905 (n13220, n_11942, n_11943);
  not g24906 (n_11944, n13220);
  and g24907 (n13221, n13217, n_11944);
  and g24908 (n13222, \a[60] , n_11941);
  and g24909 (n13223, \a[18] , n13222);
  not g24910 (n_11945, n13221);
  not g24911 (n_11946, n13223);
  and g24912 (n13224, n_11945, n_11946);
  and g24913 (n13225, n2334, n6325);
  and g24914 (n13226, n2041, n9934);
  and g24915 (n13227, n2331, n6564);
  not g24916 (n_11947, n13226);
  not g24917 (n_11948, n13227);
  and g24918 (n13228, n_11947, n_11948);
  not g24919 (n_11949, n13225);
  not g24920 (n_11950, n13228);
  and g24921 (n13229, n_11949, n_11950);
  not g24922 (n_11951, n13229);
  and g24923 (n13230, \a[51] , n_11951);
  and g24924 (n13231, \a[27] , n13230);
  and g24925 (n13232, n_11949, n_11951);
  and g24926 (n13233, \a[28] , \a[50] );
  and g24927 (n13234, \a[29] , \a[49] );
  not g24928 (n_11952, n13233);
  not g24929 (n_11953, n13234);
  and g24930 (n13235, n_11952, n_11953);
  not g24931 (n_11954, n13235);
  and g24932 (n13236, n13232, n_11954);
  not g24933 (n_11955, n13231);
  not g24934 (n_11956, n13236);
  and g24935 (n13237, n_11955, n_11956);
  not g24936 (n_11957, n13224);
  not g24937 (n_11958, n13237);
  and g24938 (n13238, n_11957, n_11958);
  not g24939 (n_11959, n13238);
  and g24940 (n13239, n_11957, n_11959);
  and g24941 (n13240, n_11958, n_11959);
  not g24942 (n_11960, n13239);
  not g24943 (n_11961, n13240);
  and g24944 (n13241, n_11960, n_11961);
  and g24945 (n13242, n1048, n9721);
  and g24946 (n13243, n993, n9909);
  and g24947 (n13244, n891, n9792);
  not g24948 (n_11962, n13243);
  not g24949 (n_11963, n13244);
  and g24950 (n13245, n_11962, n_11963);
  not g24951 (n_11964, n13242);
  not g24952 (n_11965, n13245);
  and g24953 (n13246, n_11964, n_11965);
  not g24954 (n_11966, n13246);
  and g24955 (n13247, \a[63] , n_11966);
  and g24956 (n13248, \a[15] , n13247);
  and g24957 (n13249, n_11964, n_11966);
  and g24958 (n13250, \a[16] , \a[62] );
  and g24959 (n13251, \a[17] , \a[61] );
  not g24960 (n_11967, n13250);
  not g24961 (n_11968, n13251);
  and g24962 (n13252, n_11967, n_11968);
  not g24963 (n_11969, n13252);
  and g24964 (n13253, n13249, n_11969);
  not g24965 (n_11970, n13248);
  not g24966 (n_11971, n13253);
  and g24967 (n13254, n_11970, n_11971);
  not g24968 (n_11972, n13241);
  not g24969 (n_11973, n13254);
  and g24970 (n13255, n_11972, n_11973);
  not g24971 (n_11974, n13255);
  and g24972 (n13256, n_11972, n_11974);
  and g24973 (n13257, n_11973, n_11974);
  not g24974 (n_11975, n13256);
  not g24975 (n_11976, n13257);
  and g24976 (n13258, n_11975, n_11976);
  and g24977 (n13259, \a[30] , \a[48] );
  and g24978 (n13260, \a[31] , \a[47] );
  not g24979 (n_11977, n13259);
  not g24980 (n_11978, n13260);
  and g24981 (n13261, n_11977, n_11978);
  and g24982 (n13262, n2865, n6252);
  not g24983 (n_11979, n13262);
  not g24986 (n_11980, n13261);
  not g24988 (n_11981, n13265);
  and g24989 (n13266, n_11979, n_11981);
  and g24990 (n13267, n_11980, n13266);
  and g24991 (n13268, \a[58] , n_11981);
  and g24992 (n13269, \a[20] , n13268);
  not g24993 (n_11982, n13267);
  not g24994 (n_11983, n13269);
  and g24995 (n13270, n_11982, n_11983);
  and g24996 (n13271, \a[33] , \a[45] );
  and g24997 (n13272, \a[34] , \a[44] );
  not g24998 (n_11984, n13271);
  not g24999 (n_11985, n13272);
  and g25000 (n13273, n_11984, n_11985);
  and g25001 (n13274, n4150, n5713);
  and g25002 (n13275, n4090, n7747);
  and g25003 (n13276, n3143, n5560);
  not g25004 (n_11986, n13275);
  not g25005 (n_11987, n13276);
  and g25006 (n13277, n_11986, n_11987);
  not g25007 (n_11988, n13274);
  not g25008 (n_11989, n13277);
  and g25009 (n13278, n_11988, n_11989);
  not g25010 (n_11990, n13278);
  and g25011 (n13279, n_11988, n_11990);
  not g25012 (n_11991, n13273);
  and g25013 (n13280, n_11991, n13279);
  and g25014 (n13281, n5558, n_11990);
  not g25015 (n_11992, n13280);
  not g25016 (n_11993, n13281);
  and g25017 (n13282, n_11992, n_11993);
  not g25018 (n_11994, n13270);
  not g25019 (n_11995, n13282);
  and g25020 (n13283, n_11994, n_11995);
  not g25021 (n_11996, n13283);
  and g25022 (n13284, n_11994, n_11996);
  and g25023 (n13285, n_11995, n_11996);
  not g25024 (n_11997, n13284);
  not g25025 (n_11998, n13285);
  and g25026 (n13286, n_11997, n_11998);
  and g25027 (n13287, n2115, n7421);
  and g25028 (n13288, \a[53] , \a[56] );
  and g25029 (n13289, n5327, n13288);
  and g25030 (n13290, n1904, n7699);
  not g25031 (n_11999, n13289);
  not g25032 (n_12000, n13290);
  and g25033 (n13291, n_11999, n_12000);
  not g25034 (n_12001, n13287);
  not g25035 (n_12002, n13291);
  and g25036 (n13292, n_12001, n_12002);
  not g25037 (n_12003, n13292);
  and g25038 (n13293, \a[53] , n_12003);
  and g25039 (n13294, \a[25] , n13293);
  and g25040 (n13295, \a[22] , \a[56] );
  not g25041 (n_12004, n12697);
  not g25042 (n_12005, n13295);
  and g25043 (n13296, n_12004, n_12005);
  and g25044 (n13297, n_12001, n_12003);
  not g25045 (n_12006, n13296);
  and g25046 (n13298, n_12006, n13297);
  not g25047 (n_12007, n13294);
  not g25048 (n_12008, n13298);
  and g25049 (n13299, n_12007, n_12008);
  not g25050 (n_12009, n13286);
  not g25051 (n_12010, n13299);
  and g25052 (n13300, n_12009, n_12010);
  not g25053 (n_12011, n13300);
  and g25054 (n13301, n_12009, n_12011);
  and g25055 (n13302, n_12010, n_12011);
  not g25056 (n_12012, n13301);
  not g25057 (n_12013, n13302);
  and g25058 (n13303, n_12012, n_12013);
  not g25059 (n_12014, n13258);
  and g25060 (n13304, n_12014, n13303);
  not g25061 (n_12015, n13303);
  and g25062 (n13305, n13258, n_12015);
  not g25063 (n_12016, n13304);
  not g25064 (n_12017, n13305);
  and g25065 (n13306, n_12016, n_12017);
  not g25066 (n_12018, n13210);
  not g25067 (n_12019, n13306);
  and g25068 (n13307, n_12018, n_12019);
  and g25069 (n13308, n13210, n13306);
  not g25070 (n_12020, n13307);
  not g25071 (n_12021, n13308);
  and g25072 (n13309, n_12020, n_12021);
  not g25073 (n_12022, n13209);
  and g25074 (n13310, n_12022, n13309);
  not g25075 (n_12023, n13309);
  and g25076 (n13311, n13209, n_12023);
  not g25077 (n_12024, n13310);
  not g25078 (n_12025, n13311);
  and g25079 (n13312, n_12024, n_12025);
  not g25080 (n_12026, n13312);
  and g25081 (n13313, n13208, n_12026);
  not g25082 (n_12027, n13208);
  and g25083 (n13314, n_12027, n13312);
  not g25084 (n_12028, n13313);
  not g25085 (n_12029, n13314);
  and g25086 (n13315, n_12028, n_12029);
  and g25087 (n13316, n_11775, n_11923);
  not g25088 (n_12030, n13316);
  and g25089 (n13317, n13315, n_12030);
  not g25090 (n_12031, n13315);
  and g25091 (n13318, n_12031, n13316);
  not g25092 (n_12032, n13317);
  not g25093 (n_12033, n13318);
  and g25094 (n13319, n_12032, n_12033);
  and g25095 (n13320, n_11912, n_11916);
  and g25096 (n13321, n_11841, n_11840);
  not g25097 (n_12034, n13321);
  and g25098 (n13322, n_11856, n_12034);
  and g25099 (n13323, n_11811, n_11823);
  and g25100 (n13324, n13322, n13323);
  not g25101 (n_12035, n13322);
  not g25102 (n_12036, n13323);
  and g25103 (n13325, n_12035, n_12036);
  not g25104 (n_12037, n13324);
  not g25105 (n_12038, n13325);
  and g25106 (n13326, n_12037, n_12038);
  and g25107 (n13327, n_11886, n_11898);
  not g25108 (n_12039, n13326);
  and g25109 (n13328, n_12039, n13327);
  not g25110 (n_12040, n13327);
  and g25111 (n13329, n13326, n_12040);
  not g25112 (n_12041, n13328);
  not g25113 (n_12042, n13329);
  and g25114 (n13330, n_12041, n_12042);
  and g25115 (n13331, n_11763, n_11766);
  not g25116 (n_12043, n13331);
  and g25117 (n13332, n13330, n_12043);
  not g25118 (n_12044, n13330);
  and g25119 (n13333, n_12044, n13331);
  not g25120 (n_12045, n13332);
  not g25121 (n_12046, n13333);
  and g25122 (n13334, n_12045, n_12046);
  and g25123 (n13335, n13059, n13071);
  not g25124 (n_12047, n13059);
  not g25125 (n_12048, n13071);
  and g25126 (n13336, n_12047, n_12048);
  not g25127 (n_12049, n13335);
  not g25128 (n_12050, n13336);
  and g25129 (n13337, n_12049, n_12050);
  not g25130 (n_12051, n13337);
  and g25131 (n13338, n13151, n_12051);
  not g25132 (n_12052, n13151);
  and g25133 (n13339, n_12052, n13337);
  not g25134 (n_12053, n13338);
  not g25135 (n_12054, n13339);
  and g25136 (n13340, n_12053, n_12054);
  and g25137 (n13341, n13046, n13106);
  not g25138 (n_12055, n13046);
  not g25139 (n_12056, n13106);
  and g25140 (n13342, n_12055, n_12056);
  not g25141 (n_12057, n13341);
  not g25142 (n_12058, n13342);
  and g25143 (n13343, n_12057, n_12058);
  not g25144 (n_12059, n13343);
  and g25145 (n13344, n13166, n_12059);
  not g25146 (n_12060, n13166);
  and g25147 (n13345, n_12060, n13343);
  not g25148 (n_12061, n13344);
  not g25149 (n_12062, n13345);
  and g25150 (n13346, n_12061, n_12062);
  and g25151 (n13347, n_11755, n_11759);
  not g25152 (n_12063, n13346);
  and g25153 (n13348, n_12063, n13347);
  not g25154 (n_12064, n13347);
  and g25155 (n13349, n13346, n_12064);
  not g25156 (n_12065, n13348);
  not g25157 (n_12066, n13349);
  and g25158 (n13350, n_12065, n_12066);
  and g25159 (n13351, n13340, n13350);
  not g25160 (n_12067, n13340);
  not g25161 (n_12068, n13350);
  and g25162 (n13352, n_12067, n_12068);
  not g25163 (n_12069, n13351);
  not g25164 (n_12070, n13352);
  and g25165 (n13353, n_12069, n_12070);
  and g25166 (n13354, n13334, n13353);
  not g25167 (n_12071, n13334);
  not g25168 (n_12072, n13353);
  and g25169 (n13355, n_12071, n_12072);
  not g25170 (n_12073, n13354);
  not g25171 (n_12074, n13355);
  and g25172 (n13356, n_12073, n_12074);
  not g25173 (n_12075, n13356);
  and g25174 (n13357, n13320, n_12075);
  not g25175 (n_12076, n13320);
  and g25176 (n13358, n_12076, n13356);
  not g25177 (n_12077, n13357);
  not g25178 (n_12078, n13358);
  and g25179 (n13359, n_12077, n_12078);
  and g25180 (n13360, n_11903, n_11908);
  and g25181 (n13361, n_11829, n_11861);
  not g25182 (n_12079, n13360);
  not g25183 (n_12080, n13361);
  and g25184 (n13362, n_12079, n_12080);
  not g25185 (n_12081, n13362);
  and g25186 (n13363, n_12079, n_12081);
  and g25187 (n13364, n_12080, n_12081);
  not g25188 (n_12082, n13363);
  not g25189 (n_12083, n13364);
  and g25190 (n13365, n_12082, n_12083);
  and g25191 (n13366, \a[36] , \a[42] );
  not g25192 (n_12084, n5645);
  not g25193 (n_12085, n13366);
  and g25194 (n13367, n_12084, n_12085);
  and g25195 (n13368, n3828, n5018);
  not g25196 (n_12086, n13368);
  not g25199 (n_12087, n13367);
  not g25201 (n_12088, n13371);
  and g25202 (n13372, n_12086, n_12088);
  and g25203 (n13373, n_12087, n13372);
  and g25204 (n13374, \a[55] , n_12088);
  and g25205 (n13375, \a[23] , n13374);
  not g25206 (n_12089, n13373);
  not g25207 (n_12090, n13375);
  and g25208 (n13376, n_12089, n_12090);
  and g25209 (n13377, \a[26] , \a[52] );
  and g25210 (n13378, n3803, n13377);
  and g25211 (n13379, n5946, n13377);
  and g25212 (n13380, n4565, n5413);
  not g25213 (n_12091, n13379);
  not g25214 (n_12092, n13380);
  and g25215 (n13381, n_12091, n_12092);
  not g25216 (n_12093, n13378);
  not g25217 (n_12094, n13381);
  and g25218 (n13382, n_12093, n_12094);
  not g25219 (n_12095, n13382);
  and g25220 (n13383, n5946, n_12095);
  and g25221 (n13384, n_12093, n_12095);
  not g25222 (n_12096, n3803);
  not g25223 (n_12097, n13377);
  and g25224 (n13385, n_12096, n_12097);
  not g25225 (n_12098, n13385);
  and g25226 (n13386, n13384, n_12098);
  not g25227 (n_12099, n13383);
  not g25228 (n_12100, n13386);
  and g25229 (n13387, n_12099, n_12100);
  not g25230 (n_12101, n13376);
  not g25231 (n_12102, n13387);
  and g25232 (n13388, n_12101, n_12102);
  not g25233 (n_12103, n13388);
  and g25234 (n13389, n_12101, n_12103);
  and g25235 (n13390, n_12102, n_12103);
  not g25236 (n_12104, n13389);
  not g25237 (n_12105, n13390);
  and g25238 (n13391, n_12104, n_12105);
  and g25239 (n13392, n_11747, n_11751);
  and g25240 (n13393, n13391, n13392);
  not g25241 (n_12106, n13391);
  not g25242 (n_12107, n13392);
  and g25243 (n13394, n_12106, n_12107);
  not g25244 (n_12108, n13393);
  not g25245 (n_12109, n13394);
  and g25246 (n13395, n_12108, n_12109);
  and g25247 (n13396, n13091, n13136);
  not g25248 (n_12110, n13091);
  not g25249 (n_12111, n13136);
  and g25250 (n13397, n_12110, n_12111);
  not g25251 (n_12112, n13396);
  not g25252 (n_12113, n13397);
  and g25253 (n13398, n_12112, n_12113);
  and g25254 (n13399, n_11724, n_11729);
  not g25255 (n_12114, n13398);
  and g25256 (n13400, n_12114, n13399);
  not g25257 (n_12115, n13399);
  and g25258 (n13401, n13398, n_12115);
  not g25259 (n_12116, n13400);
  not g25260 (n_12117, n13401);
  and g25261 (n13402, n_12116, n_12117);
  and g25262 (n13403, n_11735, n_11739);
  not g25263 (n_12118, n13402);
  and g25264 (n13404, n_12118, n13403);
  not g25265 (n_12119, n13403);
  and g25266 (n13405, n13402, n_12119);
  not g25267 (n_12120, n13404);
  not g25268 (n_12121, n13405);
  and g25269 (n13406, n_12120, n_12121);
  and g25270 (n13407, n13395, n13406);
  not g25271 (n_12122, n13395);
  not g25272 (n_12123, n13406);
  and g25273 (n13408, n_12122, n_12123);
  not g25274 (n_12124, n13407);
  not g25275 (n_12125, n13408);
  and g25276 (n13409, n_12124, n_12125);
  not g25277 (n_12126, n13365);
  and g25278 (n13410, n_12126, n13409);
  not g25279 (n_12127, n13410);
  and g25280 (n13411, n_12126, n_12127);
  and g25281 (n13412, n13409, n_12127);
  not g25282 (n_12128, n13411);
  not g25283 (n_12129, n13412);
  and g25284 (n13413, n_12128, n_12129);
  not g25285 (n_12130, n13413);
  and g25286 (n13414, n13359, n_12130);
  not g25287 (n_12131, n13359);
  and g25288 (n13415, n_12131, n13413);
  not g25289 (n_12132, n13415);
  and g25290 (n13416, n13319, n_12132);
  not g25291 (n_12133, n13414);
  and g25292 (n13417, n_12133, n13416);
  not g25293 (n_12134, n13417);
  and g25294 (n13418, n13319, n_12134);
  and g25295 (n13419, n_12132, n_12134);
  and g25296 (n13420, n_12133, n13419);
  not g25297 (n_12135, n13418);
  not g25298 (n_12136, n13420);
  and g25299 (n13421, n_12135, n_12136);
  not g25300 (n_12137, n13207);
  not g25301 (n_12138, n13421);
  and g25302 (n13422, n_12137, n_12138);
  and g25303 (n13423, n13207, n13421);
  not g25304 (n_12139, n13422);
  not g25305 (n_12140, n13423);
  and g25306 (n13424, n_12139, n_12140);
  not g25307 (n_12141, n13206);
  and g25308 (n13425, n_12141, n13424);
  not g25309 (n_12142, n13424);
  and g25310 (n13426, n13206, n_12142);
  not g25311 (n_12143, n13425);
  not g25312 (n_12144, n13426);
  and g25313 (\asquared[79] , n_12143, n_12144);
  and g25314 (n13428, n_12032, n_12134);
  and g25315 (n13429, n_12081, n_12127);
  and g25316 (n13430, n_12014, n_12015);
  not g25317 (n_12145, n13430);
  and g25318 (n13431, n_12020, n_12145);
  and g25319 (n13432, n13217, n13232);
  not g25320 (n_12146, n13217);
  not g25321 (n_12147, n13232);
  and g25322 (n13433, n_12146, n_12147);
  not g25323 (n_12148, n13432);
  not g25324 (n_12149, n13433);
  and g25325 (n13434, n_12148, n_12149);
  not g25326 (n_12150, n13434);
  and g25327 (n13435, n13297, n_12150);
  not g25328 (n_12151, n13297);
  and g25329 (n13436, n_12151, n13434);
  not g25330 (n_12152, n13435);
  not g25331 (n_12153, n13436);
  and g25332 (n13437, n_12152, n_12153);
  and g25333 (n13438, n_12103, n_12109);
  not g25334 (n_12154, n13437);
  and g25335 (n13439, n_12154, n13438);
  not g25336 (n_12155, n13438);
  and g25337 (n13440, n13437, n_12155);
  not g25338 (n_12156, n13439);
  not g25339 (n_12157, n13440);
  and g25340 (n13441, n_12156, n_12157);
  and g25341 (n13442, \a[34] , \a[45] );
  and g25342 (n13443, \a[35] , \a[44] );
  not g25343 (n_12158, n13442);
  not g25344 (n_12159, n13443);
  and g25345 (n13444, n_12158, n_12159);
  and g25346 (n13445, n3319, n5713);
  not g25347 (n_12160, n13445);
  not g25350 (n_12161, n13444);
  not g25352 (n_12162, n13448);
  and g25353 (n13449, n_12160, n_12162);
  and g25354 (n13450, n_12161, n13449);
  and g25355 (n13451, \a[63] , n_12162);
  and g25356 (n13452, \a[16] , n13451);
  not g25357 (n_12163, n13450);
  not g25358 (n_12164, n13452);
  and g25359 (n13453, n_12163, n_12164);
  and g25360 (n13454, \a[36] , \a[43] );
  and g25361 (n13455, \a[23] , \a[56] );
  and g25362 (n13456, \a[27] , \a[52] );
  not g25363 (n_12165, n13455);
  not g25364 (n_12166, n13456);
  and g25365 (n13457, n_12165, n_12166);
  and g25366 (n13458, \a[27] , \a[56] );
  and g25367 (n13459, n12557, n13458);
  not g25368 (n_12167, n13459);
  and g25369 (n13460, n13454, n_12167);
  not g25370 (n_12168, n13457);
  and g25371 (n13461, n_12168, n13460);
  not g25372 (n_12169, n13461);
  and g25373 (n13462, n13454, n_12169);
  and g25374 (n13463, n_12167, n_12169);
  and g25375 (n13464, n_12168, n13463);
  not g25376 (n_12170, n13462);
  not g25377 (n_12171, n13464);
  and g25378 (n13465, n_12170, n_12171);
  not g25379 (n_12172, n13453);
  not g25380 (n_12173, n13465);
  and g25381 (n13466, n_12172, n_12173);
  not g25382 (n_12174, n13466);
  and g25383 (n13467, n_12172, n_12174);
  and g25384 (n13468, n_12173, n_12174);
  not g25385 (n_12175, n13467);
  not g25386 (n_12176, n13468);
  and g25387 (n13469, n_12175, n_12176);
  and g25388 (n13470, n_12113, n_12117);
  and g25389 (n13471, n13469, n13470);
  not g25390 (n_12177, n13469);
  not g25391 (n_12178, n13470);
  and g25392 (n13472, n_12177, n_12178);
  not g25393 (n_12179, n13471);
  not g25394 (n_12180, n13472);
  and g25395 (n13473, n_12179, n_12180);
  and g25396 (n13474, n13441, n13473);
  not g25397 (n_12181, n13441);
  not g25398 (n_12182, n13473);
  and g25399 (n13475, n_12181, n_12182);
  not g25400 (n_12183, n13474);
  not g25401 (n_12184, n13475);
  and g25402 (n13476, n_12183, n_12184);
  not g25403 (n_12185, n13476);
  and g25404 (n13477, n13431, n_12185);
  not g25405 (n_12186, n13431);
  and g25406 (n13478, n_12186, n13476);
  not g25407 (n_12187, n13477);
  not g25408 (n_12188, n13478);
  and g25409 (n13479, n_12187, n_12188);
  and g25410 (n13480, n_11996, n_12011);
  and g25411 (n13481, \a[18] , \a[61] );
  not g25412 (n_12189, n13384);
  and g25413 (n13482, n_12189, n13481);
  not g25414 (n_12190, n13481);
  and g25415 (n13483, n13384, n_12190);
  not g25416 (n_12191, n13482);
  not g25417 (n_12192, n13483);
  and g25418 (n13484, n_12191, n_12192);
  not g25419 (n_12193, n13484);
  and g25420 (n13485, n13372, n_12193);
  not g25421 (n_12194, n13372);
  and g25422 (n13486, n_12194, n13484);
  not g25423 (n_12195, n13485);
  not g25424 (n_12196, n13486);
  and g25425 (n13487, n_12195, n_12196);
  and g25426 (n13488, n13249, n13266);
  not g25427 (n_12197, n13249);
  not g25428 (n_12198, n13266);
  and g25429 (n13489, n_12197, n_12198);
  not g25430 (n_12199, n13488);
  not g25431 (n_12200, n13489);
  and g25432 (n13490, n_12199, n_12200);
  not g25433 (n_12201, n13490);
  and g25434 (n13491, n13279, n_12201);
  not g25435 (n_12202, n13279);
  and g25436 (n13492, n_12202, n13490);
  not g25437 (n_12203, n13491);
  not g25438 (n_12204, n13492);
  and g25439 (n13493, n_12203, n_12204);
  and g25440 (n13494, n13487, n13493);
  not g25441 (n_12205, n13487);
  not g25442 (n_12206, n13493);
  and g25443 (n13495, n_12205, n_12206);
  not g25444 (n_12207, n13494);
  not g25445 (n_12208, n13495);
  and g25446 (n13496, n_12207, n_12208);
  not g25447 (n_12209, n13480);
  and g25448 (n13497, n_12209, n13496);
  not g25449 (n_12210, n13496);
  and g25450 (n13498, n13480, n_12210);
  not g25451 (n_12211, n13497);
  not g25452 (n_12212, n13498);
  and g25453 (n13499, n_12211, n_12212);
  and g25454 (n13500, n13479, n13499);
  not g25455 (n_12213, n13479);
  not g25456 (n_12214, n13499);
  and g25457 (n13501, n_12213, n_12214);
  not g25458 (n_12215, n13500);
  not g25459 (n_12216, n13501);
  and g25460 (n13502, n_12215, n_12216);
  not g25461 (n_12217, n13502);
  and g25462 (n13503, n13429, n_12217);
  not g25463 (n_12218, n13429);
  and g25464 (n13504, n_12218, n13502);
  not g25465 (n_12219, n13503);
  not g25466 (n_12220, n13504);
  and g25467 (n13505, n_12219, n_12220);
  and g25468 (n13506, n_12024, n_12029);
  not g25469 (n_12221, n13505);
  and g25470 (n13507, n_12221, n13506);
  not g25471 (n_12222, n13506);
  and g25472 (n13508, n13505, n_12222);
  not g25473 (n_12223, n13507);
  not g25474 (n_12224, n13508);
  and g25475 (n13509, n_12223, n_12224);
  and g25476 (n13510, n_12078, n_12133);
  and g25477 (n13511, n_12045, n_12073);
  and g25478 (n13512, n_12066, n_12069);
  and g25479 (n13513, n2463, n7699);
  and g25480 (n13514, n2301, n7697);
  and g25481 (n13515, n1904, n7701);
  not g25482 (n_12225, n13514);
  not g25483 (n_12226, n13515);
  and g25484 (n13516, n_12225, n_12226);
  not g25485 (n_12227, n13513);
  not g25486 (n_12228, n13516);
  and g25487 (n13517, n_12227, n_12228);
  not g25488 (n_12229, n13517);
  and g25489 (n13518, n_12227, n_12229);
  and g25490 (n13519, \a[25] , \a[54] );
  and g25491 (n13520, \a[26] , \a[53] );
  not g25492 (n_12230, n13519);
  not g25493 (n_12231, n13520);
  and g25494 (n13521, n_12230, n_12231);
  not g25495 (n_12232, n13521);
  and g25496 (n13522, n13518, n_12232);
  and g25497 (n13523, \a[55] , n_12229);
  and g25498 (n13524, \a[24] , n13523);
  not g25499 (n_12233, n13522);
  not g25500 (n_12234, n13524);
  and g25501 (n13525, n_12233, n_12234);
  and g25502 (n13526, \a[37] , \a[42] );
  and g25503 (n13527, n5083, n5413);
  and g25504 (n13528, n4171, n13526);
  and g25505 (n13529, n4565, n5344);
  not g25506 (n_12235, n13528);
  not g25507 (n_12236, n13529);
  and g25508 (n13530, n_12235, n_12236);
  not g25509 (n_12237, n13527);
  not g25510 (n_12238, n13530);
  and g25511 (n13531, n_12237, n_12238);
  not g25512 (n_12239, n13531);
  and g25513 (n13532, n13526, n_12239);
  and g25514 (n13533, n_12237, n_12239);
  and g25515 (n13534, \a[38] , \a[41] );
  not g25516 (n_12240, n4171);
  not g25517 (n_12241, n13534);
  and g25518 (n13535, n_12240, n_12241);
  not g25519 (n_12242, n13535);
  and g25520 (n13536, n13533, n_12242);
  not g25521 (n_12243, n13532);
  not g25522 (n_12244, n13536);
  and g25523 (n13537, n_12243, n_12244);
  not g25524 (n_12245, n13525);
  not g25525 (n_12246, n13537);
  and g25526 (n13538, n_12245, n_12246);
  not g25527 (n_12247, n13538);
  and g25528 (n13539, n_12245, n_12247);
  and g25529 (n13540, n_12246, n_12247);
  not g25530 (n_12248, n13539);
  not g25531 (n_12249, n13540);
  and g25532 (n13541, n_12248, n_12249);
  and g25533 (n13542, \a[17] , \a[62] );
  not g25534 (n_12250, \a[40] );
  not g25535 (n_12251, n13542);
  and g25536 (n13543, n_12250, n_12251);
  and g25537 (n13544, \a[40] , \a[62] );
  and g25538 (n13545, \a[17] , n13544);
  not g25539 (n_12252, n13545);
  not g25542 (n_12253, n13543);
  not g25544 (n_12254, n13548);
  and g25545 (n13549, \a[51] , n_12254);
  and g25546 (n13550, \a[28] , n13549);
  and g25547 (n13551, n_12252, n_12254);
  and g25548 (n13552, n_12253, n13551);
  not g25549 (n_12255, n13550);
  not g25550 (n_12256, n13552);
  and g25551 (n13553, n_12255, n_12256);
  not g25552 (n_12257, n13541);
  not g25553 (n_12258, n13553);
  and g25554 (n13554, n_12257, n_12258);
  not g25555 (n_12259, n13554);
  and g25556 (n13555, n_12257, n_12259);
  and g25557 (n13556, n_12258, n_12259);
  not g25558 (n_12260, n13555);
  not g25559 (n_12261, n13556);
  and g25560 (n13557, n_12260, n_12261);
  and g25561 (n13558, n1494, n8987);
  and g25562 (n13559, n1492, n10089);
  and g25563 (n13560, n1490, n9509);
  not g25564 (n_12262, n13559);
  not g25565 (n_12263, n13560);
  and g25566 (n13561, n_12262, n_12263);
  not g25567 (n_12264, n13558);
  not g25568 (n_12265, n13561);
  and g25569 (n13562, n_12264, n_12265);
  not g25570 (n_12266, n13562);
  and g25571 (n13563, n_12264, n_12266);
  and g25572 (n13564, \a[20] , \a[59] );
  and g25573 (n13565, \a[21] , \a[58] );
  not g25574 (n_12267, n13564);
  not g25575 (n_12268, n13565);
  and g25576 (n13566, n_12267, n_12268);
  not g25577 (n_12269, n13566);
  and g25578 (n13567, n13563, n_12269);
  and g25579 (n13568, \a[60] , n_12266);
  and g25580 (n13569, \a[19] , n13568);
  not g25581 (n_12270, n13567);
  not g25582 (n_12271, n13569);
  and g25583 (n13570, n_12270, n_12271);
  and g25584 (n13571, \a[22] , \a[57] );
  and g25585 (n13572, \a[29] , \a[50] );
  and g25586 (n13573, \a[30] , \a[49] );
  not g25587 (n_12272, n13572);
  not g25588 (n_12273, n13573);
  and g25589 (n13574, n_12272, n_12273);
  and g25590 (n13575, n2617, n6325);
  not g25591 (n_12274, n13575);
  and g25592 (n13576, n13571, n_12274);
  not g25593 (n_12275, n13574);
  and g25594 (n13577, n_12275, n13576);
  not g25595 (n_12276, n13577);
  and g25596 (n13578, n13571, n_12276);
  and g25597 (n13579, n_12274, n_12276);
  and g25598 (n13580, n_12275, n13579);
  not g25599 (n_12277, n13578);
  not g25600 (n_12278, n13580);
  and g25601 (n13581, n_12277, n_12278);
  not g25602 (n_12279, n13570);
  not g25603 (n_12280, n13581);
  and g25604 (n13582, n_12279, n_12280);
  not g25605 (n_12281, n13582);
  and g25606 (n13583, n_12279, n_12281);
  and g25607 (n13584, n_12280, n_12281);
  not g25608 (n_12282, n13583);
  not g25609 (n_12283, n13584);
  and g25610 (n13585, n_12282, n_12283);
  and g25611 (n13586, n3143, n5666);
  and g25612 (n13587, n2598, n8578);
  and g25613 (n13588, n3812, n6252);
  not g25614 (n_12284, n13587);
  not g25615 (n_12285, n13588);
  and g25616 (n13589, n_12284, n_12285);
  not g25617 (n_12286, n13586);
  not g25618 (n_12287, n13589);
  and g25619 (n13590, n_12286, n_12287);
  not g25620 (n_12288, n13590);
  and g25621 (n13591, \a[48] , n_12288);
  and g25622 (n13592, \a[31] , n13591);
  and g25623 (n13593, \a[32] , \a[47] );
  not g25624 (n_12289, n5896);
  not g25625 (n_12290, n13593);
  and g25626 (n13594, n_12289, n_12290);
  and g25627 (n13595, n_12286, n_12288);
  not g25628 (n_12291, n13594);
  and g25629 (n13596, n_12291, n13595);
  not g25630 (n_12292, n13592);
  not g25631 (n_12293, n13596);
  and g25632 (n13597, n_12292, n_12293);
  not g25633 (n_12294, n13585);
  not g25634 (n_12295, n13597);
  and g25635 (n13598, n_12294, n_12295);
  not g25636 (n_12296, n13598);
  and g25637 (n13599, n_12294, n_12296);
  and g25638 (n13600, n_12295, n_12296);
  not g25639 (n_12297, n13599);
  not g25640 (n_12298, n13600);
  and g25641 (n13601, n_12297, n_12298);
  and g25642 (n13602, n13557, n13601);
  not g25643 (n_12299, n13557);
  not g25644 (n_12300, n13601);
  and g25645 (n13603, n_12299, n_12300);
  not g25646 (n_12301, n13602);
  not g25647 (n_12302, n13603);
  and g25648 (n13604, n_12301, n_12302);
  not g25649 (n_12303, n13512);
  and g25650 (n13605, n_12303, n13604);
  not g25651 (n_12304, n13604);
  and g25652 (n13606, n13512, n_12304);
  not g25653 (n_12305, n13605);
  not g25654 (n_12306, n13606);
  and g25655 (n13607, n_12305, n_12306);
  not g25656 (n_12307, n13607);
  and g25657 (n13608, n13511, n_12307);
  not g25658 (n_12308, n13511);
  and g25659 (n13609, n_12308, n13607);
  not g25660 (n_12309, n13608);
  not g25661 (n_12310, n13609);
  and g25662 (n13610, n_12309, n_12310);
  and g25663 (n13611, n_12058, n_12062);
  and g25664 (n13612, n_12050, n_12054);
  and g25665 (n13613, n13611, n13612);
  not g25666 (n_12311, n13611);
  not g25667 (n_12312, n13612);
  and g25668 (n13614, n_12311, n_12312);
  not g25669 (n_12313, n13613);
  not g25670 (n_12314, n13614);
  and g25671 (n13615, n_12313, n_12314);
  and g25672 (n13616, n_11959, n_11974);
  not g25673 (n_12315, n13615);
  and g25674 (n13617, n_12315, n13616);
  not g25675 (n_12316, n13616);
  and g25676 (n13618, n13615, n_12316);
  not g25677 (n_12317, n13617);
  not g25678 (n_12318, n13618);
  and g25679 (n13619, n_12317, n_12318);
  and g25680 (n13620, n_12038, n_12042);
  not g25681 (n_12319, n13619);
  and g25682 (n13621, n_12319, n13620);
  not g25683 (n_12320, n13620);
  and g25684 (n13622, n13619, n_12320);
  not g25685 (n_12321, n13621);
  not g25686 (n_12322, n13622);
  and g25687 (n13623, n_12321, n_12322);
  and g25688 (n13624, n_12121, n_12124);
  not g25689 (n_12323, n13624);
  and g25690 (n13625, n13623, n_12323);
  not g25691 (n_12324, n13623);
  and g25692 (n13626, n_12324, n13624);
  not g25693 (n_12325, n13625);
  not g25694 (n_12326, n13626);
  and g25695 (n13627, n_12325, n_12326);
  and g25696 (n13628, n13610, n13627);
  not g25697 (n_12327, n13610);
  not g25698 (n_12328, n13627);
  and g25699 (n13629, n_12327, n_12328);
  not g25700 (n_12329, n13628);
  not g25701 (n_12330, n13629);
  and g25702 (n13630, n_12329, n_12330);
  not g25703 (n_12331, n13510);
  and g25704 (n13631, n_12331, n13630);
  not g25705 (n_12332, n13631);
  and g25706 (n13632, n13630, n_12332);
  and g25707 (n13633, n_12331, n_12332);
  not g25708 (n_12333, n13632);
  not g25709 (n_12334, n13633);
  and g25710 (n13634, n_12333, n_12334);
  not g25711 (n_12335, n13634);
  and g25712 (n13635, n13509, n_12335);
  not g25713 (n_12336, n13509);
  and g25714 (n13636, n_12336, n_12334);
  and g25715 (n13637, n_12333, n13636);
  not g25716 (n_12337, n13635);
  not g25717 (n_12338, n13637);
  and g25718 (n13638, n_12337, n_12338);
  not g25719 (n_12339, n13428);
  and g25720 (n13639, n_12339, n13638);
  not g25721 (n_12340, n13638);
  and g25722 (n13640, n13428, n_12340);
  not g25723 (n_12341, n13639);
  not g25724 (n_12342, n13640);
  and g25725 (n13641, n_12341, n_12342);
  and g25726 (n13642, n_12141, n_12140);
  not g25727 (n_12343, n13642);
  and g25728 (n13643, n_12139, n_12343);
  not g25729 (n_12344, n13641);
  and g25730 (n13644, n_12344, n13643);
  not g25731 (n_12345, n13643);
  and g25732 (n13645, n13641, n_12345);
  not g25733 (n_12346, n13644);
  not g25734 (n_12347, n13645);
  and g25735 (\asquared[80] , n_12346, n_12347);
  and g25736 (n13647, n_12342, n_12345);
  not g25737 (n_12348, n13647);
  and g25738 (n13648, n_12341, n_12348);
  and g25739 (n13649, n_12332, n_12337);
  and g25740 (n13650, n_12220, n_12224);
  and g25741 (n13651, n_12188, n_12215);
  and g25742 (n13652, n_12322, n_12325);
  and g25743 (n13653, \a[17] , \a[63] );
  and g25744 (n13654, \a[29] , \a[51] );
  not g25745 (n_12349, n13653);
  not g25746 (n_12350, n13654);
  and g25747 (n13655, n_12349, n_12350);
  and g25748 (n13656, \a[29] , \a[63] );
  and g25749 (n13657, n7772, n13656);
  not g25750 (n_12351, n13657);
  not g25753 (n_12352, n13655);
  not g25755 (n_12353, n13660);
  and g25756 (n13661, n_12351, n_12353);
  and g25757 (n13662, n_12352, n13661);
  and g25758 (n13663, \a[47] , n_12353);
  and g25759 (n13664, \a[33] , n13663);
  not g25760 (n_12354, n13662);
  not g25761 (n_12355, n13664);
  and g25762 (n13665, n_12354, n_12355);
  and g25763 (n13666, n3828, n5713);
  and g25764 (n13667, n4595, n7747);
  and g25765 (n13668, n3319, n5560);
  not g25766 (n_12356, n13667);
  not g25767 (n_12357, n13668);
  and g25768 (n13669, n_12356, n_12357);
  not g25769 (n_12358, n13666);
  not g25770 (n_12359, n13669);
  and g25771 (n13670, n_12358, n_12359);
  not g25772 (n_12360, n13670);
  and g25773 (n13671, \a[46] , n_12360);
  and g25774 (n13672, \a[34] , n13671);
  and g25775 (n13673, n_12358, n_12360);
  not g25776 (n_12361, n5848);
  not g25777 (n_12362, n5933);
  and g25778 (n13674, n_12361, n_12362);
  not g25779 (n_12363, n13674);
  and g25780 (n13675, n13673, n_12363);
  not g25781 (n_12364, n13672);
  not g25782 (n_12365, n13675);
  and g25783 (n13676, n_12364, n_12365);
  not g25784 (n_12366, n13665);
  not g25785 (n_12367, n13676);
  and g25786 (n13677, n_12366, n_12367);
  not g25787 (n_12368, n13677);
  and g25788 (n13678, n_12366, n_12368);
  and g25789 (n13679, n_12367, n_12368);
  not g25790 (n_12369, n13678);
  not g25791 (n_12370, n13679);
  and g25792 (n13680, n_12369, n_12370);
  and g25793 (n13681, n1149, n9721);
  not g25794 (n_12371, n13681);
  and g25795 (n13682, \a[61] , n_12371);
  and g25796 (n13683, \a[19] , n13682);
  and g25797 (n13684, \a[62] , n_12371);
  and g25798 (n13685, \a[18] , n13684);
  not g25799 (n_12372, n13683);
  not g25800 (n_12373, n13685);
  and g25801 (n13686, n_12372, n_12373);
  not g25802 (n_12374, n13551);
  not g25803 (n_12375, n13686);
  and g25804 (n13687, n_12374, n_12375);
  not g25805 (n_12376, n13687);
  and g25806 (n13688, n_12374, n_12376);
  and g25807 (n13689, n_12375, n_12376);
  not g25808 (n_12377, n13688);
  not g25809 (n_12378, n13689);
  and g25810 (n13690, n_12377, n_12378);
  not g25811 (n_12379, n13680);
  and g25812 (n13691, n_12379, n13690);
  not g25813 (n_12380, n13690);
  and g25814 (n13692, n13680, n_12380);
  not g25815 (n_12381, n13691);
  not g25816 (n_12382, n13692);
  and g25817 (n13693, n_12381, n_12382);
  and g25818 (n13694, n1574, n8987);
  and g25819 (n13695, n1693, n10089);
  and g25820 (n13696, n1494, n9509);
  not g25821 (n_12383, n13695);
  not g25822 (n_12384, n13696);
  and g25823 (n13697, n_12383, n_12384);
  not g25824 (n_12385, n13694);
  not g25825 (n_12386, n13697);
  and g25826 (n13698, n_12385, n_12386);
  and g25827 (n13699, \a[21] , \a[59] );
  and g25828 (n13700, \a[22] , \a[58] );
  not g25829 (n_12387, n13699);
  not g25830 (n_12388, n13700);
  and g25831 (n13701, n_12387, n_12388);
  not g25832 (n_12389, n13701);
  and g25833 (n13702, n_12385, n_12389);
  and g25834 (n13703, \a[20] , \a[60] );
  not g25835 (n_12390, n13702);
  not g25836 (n_12391, n13703);
  and g25837 (n13704, n_12390, n_12391);
  not g25838 (n_12392, n13698);
  not g25839 (n_12393, n13704);
  and g25840 (n13705, n_12392, n_12393);
  not g25841 (n_12394, n13533);
  and g25842 (n13706, n_12394, n13705);
  not g25843 (n_12395, n13705);
  and g25844 (n13707, n13533, n_12395);
  not g25845 (n_12396, n13706);
  not g25846 (n_12397, n13707);
  and g25847 (n13708, n_12396, n_12397);
  and g25848 (n13709, n3812, n6256);
  and g25849 (n13710, n2488, n5888);
  and g25850 (n13711, n2865, n6325);
  not g25851 (n_12398, n13710);
  not g25852 (n_12399, n13711);
  and g25853 (n13712, n_12398, n_12399);
  not g25854 (n_12400, n13709);
  not g25855 (n_12401, n13712);
  and g25856 (n13713, n_12400, n_12401);
  not g25857 (n_12402, n13713);
  and g25858 (n13714, \a[50] , n_12402);
  and g25859 (n13715, \a[30] , n13714);
  and g25860 (n13716, n_12400, n_12402);
  and g25861 (n13717, \a[31] , \a[49] );
  and g25862 (n13718, \a[32] , \a[48] );
  not g25863 (n_12403, n13717);
  not g25864 (n_12404, n13718);
  and g25865 (n13719, n_12403, n_12404);
  not g25866 (n_12405, n13719);
  and g25867 (n13720, n13716, n_12405);
  not g25868 (n_12406, n13715);
  not g25869 (n_12407, n13720);
  and g25870 (n13721, n_12406, n_12407);
  not g25871 (n_12408, n13721);
  and g25872 (n13722, n13708, n_12408);
  not g25873 (n_12409, n13722);
  and g25874 (n13723, n13708, n_12409);
  and g25875 (n13724, n_12408, n_12409);
  not g25876 (n_12410, n13723);
  not g25877 (n_12411, n13724);
  and g25878 (n13725, n_12410, n_12411);
  and g25879 (n13726, \a[24] , \a[56] );
  and g25880 (n13727, \a[26] , \a[54] );
  not g25881 (n_12412, n13726);
  not g25882 (n_12413, n13727);
  and g25883 (n13728, n_12412, n_12413);
  and g25884 (n13729, n2301, n7421);
  and g25885 (n13730, \a[54] , \a[57] );
  and g25886 (n13731, n2303, n13730);
  and g25887 (n13732, n1666, n8200);
  not g25888 (n_12414, n13731);
  not g25889 (n_12415, n13732);
  and g25890 (n13733, n_12414, n_12415);
  not g25891 (n_12416, n13729);
  not g25892 (n_12417, n13733);
  and g25893 (n13734, n_12416, n_12417);
  not g25894 (n_12418, n13734);
  and g25895 (n13735, n_12416, n_12418);
  not g25896 (n_12419, n13728);
  and g25897 (n13736, n_12419, n13735);
  and g25898 (n13737, \a[57] , n_12418);
  and g25899 (n13738, \a[23] , n13737);
  not g25900 (n_12420, n13736);
  not g25901 (n_12421, n13738);
  and g25902 (n13739, n_12420, n_12421);
  and g25903 (n13740, \a[25] , \a[55] );
  and g25904 (n13741, \a[37] , \a[43] );
  and g25905 (n13742, \a[38] , \a[42] );
  not g25906 (n_12422, n13741);
  not g25907 (n_12423, n13742);
  and g25908 (n13743, n_12422, n_12423);
  and g25909 (n13744, n4565, n5018);
  not g25910 (n_12424, n13744);
  and g25911 (n13745, n13740, n_12424);
  not g25912 (n_12425, n13743);
  and g25913 (n13746, n_12425, n13745);
  not g25914 (n_12426, n13746);
  and g25915 (n13747, n13740, n_12426);
  and g25916 (n13748, n_12424, n_12426);
  and g25917 (n13749, n_12425, n13748);
  not g25918 (n_12427, n13747);
  not g25919 (n_12428, n13749);
  and g25920 (n13750, n_12427, n_12428);
  not g25921 (n_12429, n13739);
  not g25922 (n_12430, n13750);
  and g25923 (n13751, n_12429, n_12430);
  not g25924 (n_12431, n13751);
  and g25925 (n13752, n_12429, n_12431);
  and g25926 (n13753, n_12430, n_12431);
  not g25927 (n_12432, n13752);
  not g25928 (n_12433, n13753);
  and g25929 (n13754, n_12432, n_12433);
  and g25930 (n13755, \a[27] , \a[53] );
  and g25931 (n13756, \a[28] , \a[52] );
  not g25932 (n_12434, n13755);
  not g25933 (n_12435, n13756);
  and g25934 (n13757, n_12434, n_12435);
  and g25935 (n13758, n2331, n7433);
  not g25936 (n_12436, n13758);
  and g25937 (n13759, n3984, n_12436);
  not g25938 (n_12437, n13757);
  and g25939 (n13760, n_12437, n13759);
  not g25940 (n_12438, n13760);
  and g25941 (n13761, n3984, n_12438);
  and g25942 (n13762, n_12436, n_12438);
  and g25943 (n13763, n_12437, n13762);
  not g25944 (n_12439, n13761);
  not g25945 (n_12440, n13763);
  and g25946 (n13764, n_12439, n_12440);
  not g25947 (n_12441, n13754);
  not g25948 (n_12442, n13764);
  and g25949 (n13765, n_12441, n_12442);
  not g25950 (n_12443, n13765);
  and g25951 (n13766, n_12441, n_12443);
  and g25952 (n13767, n_12442, n_12443);
  not g25953 (n_12444, n13766);
  not g25954 (n_12445, n13767);
  and g25955 (n13768, n_12444, n_12445);
  not g25956 (n_12446, n13725);
  and g25957 (n13769, n_12446, n13768);
  not g25958 (n_12447, n13768);
  and g25959 (n13770, n13725, n_12447);
  not g25960 (n_12448, n13769);
  not g25961 (n_12449, n13770);
  and g25962 (n13771, n_12448, n_12449);
  not g25963 (n_12450, n13693);
  not g25964 (n_12451, n13771);
  and g25965 (n13772, n_12450, n_12451);
  and g25966 (n13773, n13693, n13771);
  not g25967 (n_12452, n13772);
  not g25968 (n_12453, n13773);
  and g25969 (n13774, n_12452, n_12453);
  not g25970 (n_12454, n13652);
  and g25971 (n13775, n_12454, n13774);
  not g25972 (n_12455, n13774);
  and g25973 (n13776, n13652, n_12455);
  not g25974 (n_12456, n13775);
  not g25975 (n_12457, n13776);
  and g25976 (n13777, n_12456, n_12457);
  not g25977 (n_12458, n13651);
  and g25978 (n13778, n_12458, n13777);
  not g25979 (n_12459, n13777);
  and g25980 (n13779, n13651, n_12459);
  not g25981 (n_12460, n13778);
  not g25982 (n_12461, n13779);
  and g25983 (n13780, n_12460, n_12461);
  not g25984 (n_12462, n13780);
  and g25985 (n13781, n13650, n_12462);
  not g25986 (n_12463, n13650);
  and g25987 (n13782, n_12463, n13780);
  not g25988 (n_12464, n13781);
  not g25989 (n_12465, n13782);
  and g25990 (n13783, n_12464, n_12465);
  and g25991 (n13784, n_12310, n_12329);
  and g25992 (n13785, n_12149, n_12153);
  and g25993 (n13786, n_12200, n_12204);
  and g25994 (n13787, n13785, n13786);
  not g25995 (n_12466, n13785);
  not g25996 (n_12467, n13786);
  and g25997 (n13788, n_12466, n_12467);
  not g25998 (n_12468, n13787);
  not g25999 (n_12469, n13788);
  and g26000 (n13789, n_12468, n_12469);
  and g26001 (n13790, n_12191, n_12196);
  not g26002 (n_12470, n13789);
  and g26003 (n13791, n_12470, n13790);
  not g26004 (n_12471, n13790);
  and g26005 (n13792, n13789, n_12471);
  not g26006 (n_12472, n13791);
  not g26007 (n_12473, n13792);
  and g26008 (n13793, n_12472, n_12473);
  and g26009 (n13794, n_12157, n_12183);
  and g26010 (n13795, n_12207, n_12211);
  not g26011 (n_12474, n13794);
  not g26012 (n_12475, n13795);
  and g26013 (n13796, n_12474, n_12475);
  not g26014 (n_12476, n13796);
  and g26015 (n13797, n_12474, n_12476);
  and g26016 (n13798, n_12475, n_12476);
  not g26017 (n_12477, n13797);
  not g26018 (n_12478, n13798);
  and g26019 (n13799, n_12477, n_12478);
  not g26020 (n_12479, n13793);
  and g26021 (n13800, n_12479, n13799);
  not g26022 (n_12480, n13799);
  and g26023 (n13801, n13793, n_12480);
  not g26024 (n_12481, n13800);
  not g26025 (n_12482, n13801);
  and g26026 (n13802, n_12481, n_12482);
  and g26027 (n13803, n_12302, n_12305);
  and g26028 (n13804, n13449, n13518);
  not g26029 (n_12483, n13449);
  not g26030 (n_12484, n13518);
  and g26031 (n13805, n_12483, n_12484);
  not g26032 (n_12485, n13804);
  not g26033 (n_12486, n13805);
  and g26034 (n13806, n_12485, n_12486);
  not g26035 (n_12487, n13806);
  and g26036 (n13807, n13463, n_12487);
  not g26037 (n_12488, n13463);
  and g26038 (n13808, n_12488, n13806);
  not g26039 (n_12489, n13807);
  not g26040 (n_12490, n13808);
  and g26041 (n13809, n_12489, n_12490);
  and g26042 (n13810, n_12174, n_12180);
  not g26043 (n_12491, n13809);
  and g26044 (n13811, n_12491, n13810);
  not g26045 (n_12492, n13810);
  and g26046 (n13812, n13809, n_12492);
  not g26047 (n_12493, n13811);
  not g26048 (n_12494, n13812);
  and g26049 (n13813, n_12493, n_12494);
  and g26050 (n13814, n_12314, n_12318);
  not g26051 (n_12495, n13813);
  and g26052 (n13815, n_12495, n13814);
  not g26053 (n_12496, n13814);
  and g26054 (n13816, n13813, n_12496);
  not g26055 (n_12497, n13815);
  not g26056 (n_12498, n13816);
  and g26057 (n13817, n_12497, n_12498);
  not g26058 (n_12499, n13803);
  and g26059 (n13818, n_12499, n13817);
  not g26060 (n_12500, n13817);
  and g26061 (n13819, n13803, n_12500);
  not g26062 (n_12501, n13818);
  not g26063 (n_12502, n13819);
  and g26064 (n13820, n_12501, n_12502);
  and g26065 (n13821, n13563, n13579);
  not g26066 (n_12503, n13563);
  not g26067 (n_12504, n13579);
  and g26068 (n13822, n_12503, n_12504);
  not g26069 (n_12505, n13821);
  not g26070 (n_12506, n13822);
  and g26071 (n13823, n_12505, n_12506);
  not g26072 (n_12507, n13823);
  and g26073 (n13824, n13595, n_12507);
  not g26074 (n_12508, n13595);
  and g26075 (n13825, n_12508, n13823);
  not g26076 (n_12509, n13824);
  not g26077 (n_12510, n13825);
  and g26078 (n13826, n_12509, n_12510);
  and g26079 (n13827, n_12247, n_12259);
  and g26080 (n13828, n_12281, n_12296);
  and g26081 (n13829, n13827, n13828);
  not g26082 (n_12511, n13827);
  not g26083 (n_12512, n13828);
  and g26084 (n13830, n_12511, n_12512);
  not g26085 (n_12513, n13829);
  not g26086 (n_12514, n13830);
  and g26087 (n13831, n_12513, n_12514);
  and g26088 (n13832, n13826, n13831);
  not g26089 (n_12515, n13826);
  not g26090 (n_12516, n13831);
  and g26091 (n13833, n_12515, n_12516);
  not g26092 (n_12517, n13832);
  not g26093 (n_12518, n13833);
  and g26094 (n13834, n_12517, n_12518);
  and g26095 (n13835, n13820, n13834);
  not g26096 (n_12519, n13820);
  not g26097 (n_12520, n13834);
  and g26098 (n13836, n_12519, n_12520);
  not g26099 (n_12521, n13835);
  not g26100 (n_12522, n13836);
  and g26101 (n13837, n_12521, n_12522);
  and g26102 (n13838, n13802, n13837);
  not g26103 (n_12523, n13838);
  and g26104 (n13839, n13837, n_12523);
  and g26105 (n13840, n13802, n_12523);
  not g26106 (n_12524, n13839);
  not g26107 (n_12525, n13840);
  and g26108 (n13841, n_12524, n_12525);
  not g26109 (n_12526, n13784);
  not g26110 (n_12527, n13841);
  and g26111 (n13842, n_12526, n_12527);
  and g26112 (n13843, n13784, n_12525);
  and g26113 (n13844, n_12524, n13843);
  not g26114 (n_12528, n13842);
  not g26115 (n_12529, n13844);
  and g26116 (n13845, n_12528, n_12529);
  and g26117 (n13846, n13783, n13845);
  not g26118 (n_12530, n13783);
  not g26119 (n_12531, n13845);
  and g26120 (n13847, n_12530, n_12531);
  not g26121 (n_12532, n13846);
  not g26122 (n_12533, n13847);
  and g26123 (n13848, n_12532, n_12533);
  not g26124 (n_12534, n13848);
  and g26125 (n13849, n13649, n_12534);
  not g26126 (n_12535, n13649);
  and g26127 (n13850, n_12535, n13848);
  not g26128 (n_12536, n13849);
  not g26129 (n_12537, n13850);
  and g26130 (n13851, n_12536, n_12537);
  not g26131 (n_12538, n13851);
  and g26132 (n13852, n13648, n_12538);
  not g26133 (n_12539, n13648);
  and g26134 (n13853, n_12539, n_12536);
  and g26135 (n13854, n_12537, n13853);
  not g26136 (n_12540, n13852);
  not g26137 (n_12541, n13854);
  and g26138 (\asquared[81] , n_12540, n_12541);
  not g26139 (n_12542, n13853);
  and g26140 (n13856, n_12537, n_12542);
  and g26141 (n13857, n_12523, n_12528);
  and g26142 (n13858, n_12501, n_12521);
  and g26143 (n13859, n_12476, n_12482);
  and g26144 (n13860, \a[41] , \a[62] );
  and g26145 (n13861, \a[19] , n13860);
  not g26146 (n_12543, n13861);
  and g26147 (n13862, n5413, n_12543);
  not g26148 (n_12544, n13862);
  and g26149 (n13863, n_12543, n_12544);
  and g26150 (n13864, \a[19] , \a[62] );
  not g26151 (n_12545, \a[41] );
  not g26152 (n_12546, n13864);
  and g26153 (n13865, n_12545, n_12546);
  not g26154 (n_12547, n13865);
  and g26155 (n13866, n13863, n_12547);
  and g26156 (n13867, n5413, n_12544);
  not g26157 (n_12548, n13866);
  not g26158 (n_12549, n13867);
  and g26159 (n13868, n_12548, n_12549);
  and g26160 (n13869, n1547, n7942);
  and g26161 (n13870, \a[56] , \a[59] );
  and g26162 (n13871, n5327, n13870);
  and g26163 (n13872, n1919, n8987);
  not g26164 (n_12550, n13871);
  not g26165 (n_12551, n13872);
  and g26166 (n13873, n_12550, n_12551);
  not g26167 (n_12552, n13869);
  not g26168 (n_12553, n13873);
  and g26169 (n13874, n_12552, n_12553);
  not g26170 (n_12554, n13874);
  and g26171 (n13875, \a[59] , n_12554);
  and g26172 (n13876, \a[22] , n13875);
  and g26173 (n13877, n_12552, n_12554);
  and g26174 (n13878, \a[23] , \a[58] );
  not g26175 (n_12555, n12356);
  not g26176 (n_12556, n13878);
  and g26177 (n13879, n_12555, n_12556);
  not g26178 (n_12557, n13879);
  and g26179 (n13880, n13877, n_12557);
  not g26180 (n_12558, n13876);
  not g26181 (n_12559, n13880);
  and g26182 (n13881, n_12558, n_12559);
  not g26183 (n_12560, n13868);
  not g26184 (n_12561, n13881);
  and g26185 (n13882, n_12560, n_12561);
  not g26186 (n_12562, n13882);
  and g26187 (n13883, n_12560, n_12562);
  and g26188 (n13884, n_12561, n_12562);
  not g26189 (n_12563, n13883);
  not g26190 (n_12564, n13884);
  and g26191 (n13885, n_12563, n_12564);
  and g26192 (n13886, \a[33] , \a[48] );
  and g26193 (n13887, \a[34] , \a[47] );
  not g26194 (n_12565, n13886);
  not g26195 (n_12566, n13887);
  and g26196 (n13888, n_12565, n_12566);
  and g26197 (n13889, n4150, n6252);
  not g26198 (n_12567, n13889);
  and g26199 (n13890, n10301, n_12567);
  not g26200 (n_12568, n13888);
  and g26201 (n13891, n_12568, n13890);
  not g26202 (n_12569, n13891);
  and g26203 (n13892, n10301, n_12569);
  and g26204 (n13893, n_12567, n_12569);
  and g26205 (n13894, n_12568, n13893);
  not g26206 (n_12570, n13892);
  not g26207 (n_12571, n13894);
  and g26208 (n13895, n_12570, n_12571);
  not g26209 (n_12572, n13885);
  not g26210 (n_12573, n13895);
  and g26211 (n13896, n_12572, n_12573);
  not g26212 (n_12574, n13896);
  and g26213 (n13897, n_12572, n_12574);
  and g26214 (n13898, n_12573, n_12574);
  not g26215 (n_12575, n13897);
  not g26216 (n_12576, n13898);
  and g26217 (n13899, n_12575, n_12576);
  and g26218 (n13900, n_12469, n_12473);
  and g26219 (n13901, n13899, n13900);
  not g26220 (n_12577, n13899);
  not g26221 (n_12578, n13900);
  and g26222 (n13902, n_12577, n_12578);
  not g26223 (n_12579, n13901);
  not g26224 (n_12580, n13902);
  and g26225 (n13903, n_12579, n_12580);
  and g26226 (n13904, n1494, n9512);
  and g26227 (n13905, n3648, n11634);
  and g26228 (n13906, n1331, n9909);
  not g26229 (n_12581, n13905);
  not g26230 (n_12582, n13906);
  and g26231 (n13907, n_12581, n_12582);
  not g26232 (n_12583, n13904);
  not g26233 (n_12584, n13907);
  and g26234 (n13908, n_12583, n_12584);
  not g26235 (n_12585, n13908);
  and g26236 (n13909, n_12583, n_12585);
  and g26237 (n13910, \a[20] , \a[61] );
  and g26238 (n13911, \a[21] , \a[60] );
  not g26239 (n_12586, n13910);
  not g26240 (n_12587, n13911);
  and g26241 (n13912, n_12586, n_12587);
  not g26242 (n_12588, n13912);
  and g26243 (n13913, n13909, n_12588);
  and g26244 (n13914, \a[63] , n_12585);
  and g26245 (n13915, \a[18] , n13914);
  not g26246 (n_12589, n13913);
  not g26247 (n_12590, n13915);
  and g26248 (n13916, n_12589, n_12590);
  and g26249 (n13917, \a[35] , \a[46] );
  and g26250 (n13918, n3687, n5713);
  and g26251 (n13919, n3828, n5560);
  and g26252 (n13920, \a[37] , \a[44] );
  and g26253 (n13921, n13917, n13920);
  not g26254 (n_12591, n13919);
  not g26255 (n_12592, n13921);
  and g26256 (n13922, n_12591, n_12592);
  not g26257 (n_12593, n13918);
  not g26258 (n_12594, n13922);
  and g26259 (n13923, n_12593, n_12594);
  not g26260 (n_12595, n13923);
  and g26261 (n13924, n13917, n_12595);
  and g26262 (n13925, \a[36] , \a[45] );
  not g26263 (n_12596, n13920);
  not g26264 (n_12597, n13925);
  and g26265 (n13926, n_12596, n_12597);
  and g26266 (n13927, n_12593, n_12595);
  not g26267 (n_12598, n13926);
  and g26268 (n13928, n_12598, n13927);
  not g26269 (n_12599, n13924);
  not g26270 (n_12600, n13928);
  and g26271 (n13929, n_12599, n_12600);
  not g26272 (n_12601, n13916);
  not g26273 (n_12602, n13929);
  and g26274 (n13930, n_12601, n_12602);
  not g26275 (n_12603, n13930);
  and g26276 (n13931, n_12601, n_12603);
  and g26277 (n13932, n_12602, n_12603);
  not g26278 (n_12604, n13931);
  not g26279 (n_12605, n13932);
  and g26280 (n13933, n_12604, n_12605);
  and g26281 (n13934, \a[29] , n13377);
  and g26282 (n13935, \a[53] , n2800);
  not g26283 (n_12606, n13934);
  not g26284 (n_12607, n13935);
  and g26285 (n13936, n_12606, n_12607);
  and g26286 (n13937, n2334, n7433);
  not g26287 (n_12608, n13937);
  and g26288 (n13938, \a[55] , n_12608);
  not g26289 (n_12609, n13936);
  and g26290 (n13939, n_12609, n13938);
  not g26291 (n_12610, n13939);
  and g26292 (n13940, \a[55] , n_12610);
  and g26293 (n13941, \a[26] , n13940);
  and g26294 (n13942, \a[28] , \a[53] );
  and g26295 (n13943, \a[29] , \a[52] );
  not g26296 (n_12611, n13942);
  not g26297 (n_12612, n13943);
  and g26298 (n13944, n_12611, n_12612);
  and g26299 (n13945, n_12608, n_12610);
  not g26300 (n_12613, n13944);
  and g26301 (n13946, n_12613, n13945);
  not g26302 (n_12614, n13941);
  not g26303 (n_12615, n13946);
  and g26304 (n13947, n_12614, n_12615);
  not g26305 (n_12616, n13933);
  not g26306 (n_12617, n13947);
  and g26307 (n13948, n_12616, n_12617);
  not g26308 (n_12618, n13948);
  and g26309 (n13949, n_12616, n_12618);
  and g26310 (n13950, n_12617, n_12618);
  not g26311 (n_12619, n13949);
  not g26312 (n_12620, n13950);
  and g26313 (n13951, n_12619, n_12620);
  not g26314 (n_12621, n13903);
  and g26315 (n13952, n_12621, n13951);
  not g26316 (n_12622, n13951);
  and g26317 (n13953, n13903, n_12622);
  not g26318 (n_12623, n13952);
  not g26319 (n_12624, n13953);
  and g26320 (n13954, n_12623, n_12624);
  not g26321 (n_12625, n13859);
  and g26322 (n13955, n_12625, n13954);
  not g26323 (n_12626, n13955);
  and g26324 (n13956, n_12625, n_12626);
  and g26325 (n13957, n13954, n_12626);
  not g26326 (n_12627, n13956);
  not g26327 (n_12628, n13957);
  and g26328 (n13958, n_12627, n_12628);
  not g26329 (n_12629, n13858);
  not g26330 (n_12630, n13958);
  and g26331 (n13959, n_12629, n_12630);
  not g26332 (n_12631, n13959);
  and g26333 (n13960, n_12629, n_12631);
  and g26334 (n13961, n_12630, n_12631);
  not g26335 (n_12632, n13960);
  not g26336 (n_12633, n13961);
  and g26337 (n13962, n_12632, n_12633);
  not g26338 (n_12634, n13857);
  not g26339 (n_12635, n13962);
  and g26340 (n13963, n_12634, n_12635);
  not g26341 (n_12636, n13963);
  and g26342 (n13964, n_12634, n_12636);
  and g26343 (n13965, n_12635, n_12636);
  not g26344 (n_12637, n13964);
  not g26345 (n_12638, n13965);
  and g26346 (n13966, n_12637, n_12638);
  and g26347 (n13967, n_12456, n_12460);
  and g26348 (n13968, n_12506, n_12510);
  and g26349 (n13969, \a[27] , \a[54] );
  and g26350 (n13970, \a[38] , \a[43] );
  and g26351 (n13971, \a[39] , \a[42] );
  not g26352 (n_12639, n13970);
  not g26353 (n_12640, n13971);
  and g26354 (n13972, n_12639, n_12640);
  and g26355 (n13973, n5018, n5083);
  not g26356 (n_12641, n13973);
  and g26357 (n13974, n13969, n_12641);
  not g26358 (n_12642, n13972);
  and g26359 (n13975, n_12642, n13974);
  not g26360 (n_12643, n13975);
  and g26361 (n13976, n13969, n_12643);
  and g26362 (n13977, n_12641, n_12643);
  and g26363 (n13978, n_12642, n13977);
  not g26364 (n_12644, n13976);
  not g26365 (n_12645, n13978);
  and g26366 (n13979, n_12644, n_12645);
  not g26367 (n_12646, n13968);
  not g26368 (n_12647, n13979);
  and g26369 (n13980, n_12646, n_12647);
  not g26370 (n_12648, n13980);
  and g26371 (n13981, n_12646, n_12648);
  and g26372 (n13982, n_12647, n_12648);
  not g26373 (n_12649, n13981);
  not g26374 (n_12650, n13982);
  and g26375 (n13983, n_12649, n_12650);
  and g26376 (n13984, n_12486, n_12490);
  and g26377 (n13985, n13983, n13984);
  not g26378 (n_12651, n13983);
  not g26379 (n_12652, n13984);
  and g26380 (n13986, n_12651, n_12652);
  not g26381 (n_12653, n13985);
  not g26382 (n_12654, n13986);
  and g26383 (n13987, n_12653, n_12654);
  and g26384 (n13988, n_12494, n_12498);
  and g26385 (n13989, n_12514, n_12517);
  not g26386 (n_12655, n13988);
  not g26387 (n_12656, n13989);
  and g26388 (n13990, n_12655, n_12656);
  not g26389 (n_12657, n13990);
  and g26390 (n13991, n_12655, n_12657);
  and g26391 (n13992, n_12656, n_12657);
  not g26392 (n_12658, n13991);
  not g26393 (n_12659, n13992);
  and g26394 (n13993, n_12658, n_12659);
  not g26395 (n_12660, n13993);
  and g26396 (n13994, n13987, n_12660);
  not g26397 (n_12661, n13987);
  and g26398 (n13995, n_12661, n13993);
  not g26399 (n_12662, n13967);
  not g26400 (n_12663, n13995);
  and g26401 (n13996, n_12662, n_12663);
  not g26402 (n_12664, n13994);
  and g26403 (n13997, n_12664, n13996);
  not g26404 (n_12665, n13997);
  and g26405 (n13998, n_12662, n_12665);
  and g26406 (n13999, n_12663, n_12665);
  and g26407 (n14000, n_12664, n13999);
  not g26408 (n_12666, n13998);
  not g26409 (n_12667, n14000);
  and g26410 (n14001, n_12666, n_12667);
  and g26411 (n14002, n_12371, n_12376);
  and g26412 (n14003, n13673, n14002);
  not g26413 (n_12668, n13673);
  not g26414 (n_12669, n14002);
  and g26415 (n14004, n_12668, n_12669);
  not g26416 (n_12670, n14003);
  not g26417 (n_12671, n14004);
  and g26418 (n14005, n_12670, n_12671);
  and g26419 (n14006, n3812, n6325);
  and g26420 (n14007, n2488, n9934);
  and g26421 (n14008, n2865, n6564);
  not g26422 (n_12672, n14007);
  not g26423 (n_12673, n14008);
  and g26424 (n14009, n_12672, n_12673);
  not g26425 (n_12674, n14006);
  not g26426 (n_12675, n14009);
  and g26427 (n14010, n_12674, n_12675);
  not g26428 (n_12676, n14010);
  and g26429 (n14011, \a[51] , n_12676);
  and g26430 (n14012, \a[30] , n14011);
  and g26431 (n14013, n_12674, n_12676);
  and g26432 (n14014, \a[31] , \a[50] );
  and g26433 (n14015, \a[32] , \a[49] );
  not g26434 (n_12677, n14014);
  not g26435 (n_12678, n14015);
  and g26436 (n14016, n_12677, n_12678);
  not g26437 (n_12679, n14016);
  and g26438 (n14017, n14013, n_12679);
  not g26439 (n_12680, n14012);
  not g26440 (n_12681, n14017);
  and g26441 (n14018, n_12680, n_12681);
  not g26442 (n_12682, n14018);
  and g26443 (n14019, n14005, n_12682);
  not g26444 (n_12683, n14019);
  and g26445 (n14020, n14005, n_12683);
  and g26446 (n14021, n_12682, n_12683);
  not g26447 (n_12684, n14020);
  not g26448 (n_12685, n14021);
  and g26449 (n14022, n_12684, n_12685);
  and g26450 (n14023, n13661, n13716);
  not g26451 (n_12686, n13661);
  not g26452 (n_12687, n13716);
  and g26453 (n14024, n_12686, n_12687);
  not g26454 (n_12688, n14023);
  not g26455 (n_12689, n14024);
  and g26456 (n14025, n_12688, n_12689);
  and g26457 (n14026, n_12385, n_12392);
  not g26458 (n_12690, n14025);
  and g26459 (n14027, n_12690, n14026);
  not g26460 (n_12691, n14026);
  and g26461 (n14028, n14025, n_12691);
  not g26462 (n_12692, n14027);
  not g26463 (n_12693, n14028);
  and g26464 (n14029, n_12692, n_12693);
  and g26465 (n14030, n_12379, n_12380);
  not g26466 (n_12694, n14030);
  and g26467 (n14031, n_12368, n_12694);
  not g26468 (n_12695, n14031);
  and g26469 (n14032, n14029, n_12695);
  not g26470 (n_12696, n14029);
  and g26471 (n14033, n_12696, n14031);
  not g26472 (n_12697, n14032);
  not g26473 (n_12698, n14033);
  and g26474 (n14034, n_12697, n_12698);
  and g26475 (n14035, n14022, n14034);
  not g26476 (n_12699, n14022);
  not g26477 (n_12700, n14034);
  and g26478 (n14036, n_12699, n_12700);
  not g26479 (n_12701, n14035);
  not g26480 (n_12702, n14036);
  and g26481 (n14037, n_12701, n_12702);
  and g26482 (n14038, n_12446, n_12447);
  not g26483 (n_12703, n14038);
  and g26484 (n14039, n_12452, n_12703);
  and g26485 (n14040, n14037, n14039);
  not g26486 (n_12704, n14037);
  not g26487 (n_12705, n14039);
  and g26488 (n14041, n_12704, n_12705);
  not g26489 (n_12706, n14040);
  not g26490 (n_12707, n14041);
  and g26491 (n14042, n_12706, n_12707);
  and g26492 (n14043, n13748, n13762);
  not g26493 (n_12708, n13748);
  not g26494 (n_12709, n13762);
  and g26495 (n14044, n_12708, n_12709);
  not g26496 (n_12710, n14043);
  not g26497 (n_12711, n14044);
  and g26498 (n14045, n_12710, n_12711);
  not g26499 (n_12712, n14045);
  and g26500 (n14046, n13735, n_12712);
  not g26501 (n_12713, n13735);
  and g26502 (n14047, n_12713, n14045);
  not g26503 (n_12714, n14046);
  not g26504 (n_12715, n14047);
  and g26505 (n14048, n_12714, n_12715);
  and g26506 (n14049, n_12431, n_12443);
  and g26507 (n14050, n_12396, n_12409);
  and g26508 (n14051, n14049, n14050);
  not g26509 (n_12716, n14049);
  not g26510 (n_12717, n14050);
  and g26511 (n14052, n_12716, n_12717);
  not g26512 (n_12718, n14051);
  not g26513 (n_12719, n14052);
  and g26514 (n14053, n_12718, n_12719);
  and g26515 (n14054, n14048, n14053);
  not g26516 (n_12720, n14048);
  not g26517 (n_12721, n14053);
  and g26518 (n14055, n_12720, n_12721);
  not g26519 (n_12722, n14054);
  not g26520 (n_12723, n14055);
  and g26521 (n14056, n_12722, n_12723);
  and g26522 (n14057, n14042, n14056);
  not g26523 (n_12724, n14042);
  not g26524 (n_12725, n14056);
  and g26525 (n14058, n_12724, n_12725);
  not g26526 (n_12726, n14057);
  not g26527 (n_12727, n14058);
  and g26528 (n14059, n_12726, n_12727);
  not g26529 (n_12728, n14001);
  not g26530 (n_12729, n14059);
  and g26531 (n14060, n_12728, n_12729);
  and g26532 (n14061, n14001, n14059);
  not g26533 (n_12730, n14060);
  not g26534 (n_12731, n14061);
  and g26535 (n14062, n_12730, n_12731);
  not g26536 (n_12732, n13966);
  not g26537 (n_12733, n14062);
  and g26538 (n14063, n_12732, n_12733);
  not g26539 (n_12734, n14063);
  and g26540 (n14064, n_12732, n_12734);
  and g26541 (n14065, n_12733, n_12734);
  not g26542 (n_12735, n14064);
  not g26543 (n_12736, n14065);
  and g26544 (n14066, n_12735, n_12736);
  and g26545 (n14067, n_12465, n_12532);
  not g26546 (n_12737, n14066);
  not g26547 (n_12738, n14067);
  and g26548 (n14068, n_12737, n_12738);
  and g26549 (n14069, n14066, n14067);
  not g26550 (n_12739, n14068);
  not g26551 (n_12740, n14069);
  and g26552 (n14070, n_12739, n_12740);
  not g26553 (n_12741, n13856);
  not g26554 (n_12742, n14070);
  and g26555 (n14071, n_12741, n_12742);
  and g26556 (n14072, n13856, n14070);
  or g26557 (\asquared[82] , n14071, n14072);
  and g26558 (n14074, n_12741, n_12740);
  not g26559 (n_12743, n14074);
  and g26560 (n14075, n_12739, n_12743);
  and g26561 (n14076, n_12636, n_12734);
  and g26562 (n14077, n_12728, n14059);
  not g26563 (n_12744, n14077);
  and g26564 (n14078, n_12665, n_12744);
  and g26565 (n14079, n_12707, n_12726);
  and g26566 (n14080, n_12657, n_12664);
  and g26567 (n14081, \a[51] , \a[62] );
  and g26568 (n14082, n6098, n14081);
  and g26569 (n14083, n1494, n9721);
  not g26570 (n_12745, n14082);
  not g26571 (n_12746, n14083);
  and g26572 (n14084, n_12745, n_12746);
  and g26573 (n14085, \a[31] , \a[51] );
  and g26574 (n14086, \a[21] , \a[61] );
  and g26575 (n14087, n14085, n14086);
  not g26576 (n_12747, n14084);
  not g26577 (n_12748, n14087);
  and g26578 (n14088, n_12747, n_12748);
  not g26579 (n_12749, n14088);
  and g26580 (n14089, n_12748, n_12749);
  not g26581 (n_12750, n14085);
  not g26582 (n_12751, n14086);
  and g26583 (n14090, n_12750, n_12751);
  not g26584 (n_12752, n14090);
  and g26585 (n14091, n14089, n_12752);
  and g26586 (n14092, \a[62] , n_12749);
  and g26587 (n14093, \a[20] , n14092);
  not g26588 (n_12753, n14091);
  not g26589 (n_12754, n14093);
  and g26590 (n14094, n_12753, n_12754);
  and g26591 (n14095, n4150, n6256);
  and g26592 (n14096, n4090, n5888);
  and g26593 (n14097, n3143, n6325);
  not g26594 (n_12755, n14096);
  not g26595 (n_12756, n14097);
  and g26596 (n14098, n_12755, n_12756);
  not g26597 (n_12757, n14095);
  not g26598 (n_12758, n14098);
  and g26599 (n14099, n_12757, n_12758);
  not g26600 (n_12759, n14099);
  and g26601 (n14100, \a[50] , n_12759);
  and g26602 (n14101, \a[32] , n14100);
  and g26603 (n14102, n_12757, n_12759);
  and g26604 (n14103, \a[33] , \a[49] );
  and g26605 (n14104, \a[34] , \a[48] );
  not g26606 (n_12760, n14103);
  not g26607 (n_12761, n14104);
  and g26608 (n14105, n_12760, n_12761);
  not g26609 (n_12762, n14105);
  and g26610 (n14106, n14102, n_12762);
  not g26611 (n_12763, n14101);
  not g26612 (n_12764, n14106);
  and g26613 (n14107, n_12763, n_12764);
  not g26614 (n_12765, n14094);
  not g26615 (n_12766, n14107);
  and g26616 (n14108, n_12765, n_12766);
  not g26617 (n_12767, n14108);
  and g26618 (n14109, n_12765, n_12767);
  and g26619 (n14110, n_12766, n_12767);
  not g26620 (n_12768, n14109);
  not g26621 (n_12769, n14110);
  and g26622 (n14111, n_12768, n_12769);
  and g26623 (n14112, n1666, n8987);
  and g26624 (n14113, n2115, n10089);
  and g26625 (n14114, n1919, n9509);
  not g26626 (n_12770, n14113);
  not g26627 (n_12771, n14114);
  and g26628 (n14115, n_12770, n_12771);
  not g26629 (n_12772, n14112);
  not g26630 (n_12773, n14115);
  and g26631 (n14116, n_12772, n_12773);
  not g26632 (n_12774, n14116);
  and g26633 (n14117, \a[60] , n_12774);
  and g26634 (n14118, \a[22] , n14117);
  and g26635 (n14119, n_12772, n_12774);
  and g26636 (n14120, \a[23] , \a[59] );
  not g26637 (n_12775, n11415);
  not g26638 (n_12776, n14120);
  and g26639 (n14121, n_12775, n_12776);
  not g26640 (n_12777, n14121);
  and g26641 (n14122, n14119, n_12777);
  not g26642 (n_12778, n14118);
  not g26643 (n_12779, n14122);
  and g26644 (n14123, n_12778, n_12779);
  not g26645 (n_12780, n14111);
  not g26646 (n_12781, n14123);
  and g26647 (n14124, n_12780, n_12781);
  not g26648 (n_12782, n14124);
  and g26649 (n14125, n_12780, n_12782);
  and g26650 (n14126, n_12781, n_12782);
  not g26651 (n_12783, n14125);
  not g26652 (n_12784, n14126);
  and g26653 (n14127, n_12783, n_12784);
  and g26654 (n14128, n_12648, n_12654);
  and g26655 (n14129, n14127, n14128);
  not g26656 (n_12785, n14127);
  not g26657 (n_12786, n14128);
  and g26658 (n14130, n_12785, n_12786);
  not g26659 (n_12787, n14129);
  not g26660 (n_12788, n14130);
  and g26661 (n14131, n_12787, n_12788);
  and g26662 (n14132, \a[38] , \a[44] );
  and g26663 (n14133, \a[39] , \a[43] );
  not g26664 (n_12789, n14132);
  not g26665 (n_12790, n14133);
  and g26666 (n14134, n_12789, n_12790);
  and g26667 (n14135, n5083, n5296);
  not g26668 (n_12791, n14135);
  not g26671 (n_12792, n14134);
  not g26673 (n_12793, n14138);
  and g26674 (n14139, n_12791, n_12793);
  and g26675 (n14140, n_12792, n14139);
  and g26676 (n14141, \a[56] , n_12793);
  and g26677 (n14142, \a[26] , n14141);
  not g26678 (n_12794, n14140);
  not g26679 (n_12795, n14142);
  and g26680 (n14143, n_12794, n_12795);
  and g26681 (n14144, \a[29] , \a[53] );
  and g26682 (n14145, \a[30] , \a[52] );
  not g26683 (n_12796, n14144);
  not g26684 (n_12797, n14145);
  and g26685 (n14146, n_12796, n_12797);
  and g26686 (n14147, n2617, n7433);
  not g26687 (n_12798, n14147);
  and g26688 (n14148, n6453, n_12798);
  not g26689 (n_12799, n14146);
  and g26690 (n14149, n_12799, n14148);
  not g26691 (n_12800, n14149);
  and g26692 (n14150, n6453, n_12800);
  and g26693 (n14151, n_12798, n_12800);
  and g26694 (n14152, n_12799, n14151);
  not g26695 (n_12801, n14150);
  not g26696 (n_12802, n14152);
  and g26697 (n14153, n_12801, n_12802);
  not g26698 (n_12803, n14143);
  not g26699 (n_12804, n14153);
  and g26700 (n14154, n_12803, n_12804);
  not g26701 (n_12805, n14154);
  and g26702 (n14155, n_12803, n_12805);
  and g26703 (n14156, n_12804, n_12805);
  not g26704 (n_12806, n14155);
  not g26705 (n_12807, n14156);
  and g26706 (n14157, n_12806, n_12807);
  and g26707 (n14158, n3687, n5560);
  and g26708 (n14159, \a[37] , \a[47] );
  and g26709 (n14160, n5848, n14159);
  and g26710 (n14161, n3828, n5666);
  not g26711 (n_12808, n14160);
  not g26712 (n_12809, n14161);
  and g26713 (n14162, n_12808, n_12809);
  not g26714 (n_12810, n14158);
  not g26715 (n_12811, n14162);
  and g26716 (n14163, n_12810, n_12811);
  not g26717 (n_12812, n14163);
  and g26718 (n14164, \a[47] , n_12812);
  and g26719 (n14165, \a[35] , n14164);
  and g26720 (n14166, n_12810, n_12812);
  not g26721 (n_12813, n6146);
  not g26722 (n_12814, n6437);
  and g26723 (n14167, n_12813, n_12814);
  not g26724 (n_12815, n14167);
  and g26725 (n14168, n14166, n_12815);
  not g26726 (n_12816, n14165);
  not g26727 (n_12817, n14168);
  and g26728 (n14169, n_12816, n_12817);
  not g26729 (n_12818, n14157);
  not g26730 (n_12819, n14169);
  and g26731 (n14170, n_12818, n_12819);
  not g26732 (n_12820, n14170);
  and g26733 (n14171, n_12818, n_12820);
  and g26734 (n14172, n_12819, n_12820);
  not g26735 (n_12821, n14171);
  not g26736 (n_12822, n14172);
  and g26737 (n14173, n_12821, n_12822);
  not g26738 (n_12823, n14131);
  and g26739 (n14174, n_12823, n14173);
  not g26740 (n_12824, n14173);
  and g26741 (n14175, n14131, n_12824);
  not g26742 (n_12825, n14174);
  not g26743 (n_12826, n14175);
  and g26744 (n14176, n_12825, n_12826);
  not g26745 (n_12827, n14080);
  and g26746 (n14177, n_12827, n14176);
  not g26747 (n_12828, n14177);
  and g26748 (n14178, n_12827, n_12828);
  and g26749 (n14179, n14176, n_12828);
  not g26750 (n_12829, n14178);
  not g26751 (n_12830, n14179);
  and g26752 (n14180, n_12829, n_12830);
  not g26753 (n_12831, n14079);
  not g26754 (n_12832, n14180);
  and g26755 (n14181, n_12831, n_12832);
  not g26756 (n_12833, n14181);
  and g26757 (n14182, n_12831, n_12833);
  and g26758 (n14183, n_12832, n_12833);
  not g26759 (n_12834, n14182);
  not g26760 (n_12835, n14183);
  and g26761 (n14184, n_12834, n_12835);
  not g26762 (n_12836, n14078);
  not g26763 (n_12837, n14184);
  and g26764 (n14185, n_12836, n_12837);
  not g26765 (n_12838, n14185);
  and g26766 (n14186, n_12836, n_12838);
  and g26767 (n14187, n_12837, n_12838);
  not g26768 (n_12839, n14186);
  not g26769 (n_12840, n14187);
  and g26770 (n14188, n_12839, n_12840);
  and g26771 (n14189, n_12626, n_12631);
  and g26772 (n14190, n_12689, n_12693);
  and g26773 (n14191, n2633, n11718);
  and g26774 (n14192, n2331, n7701);
  and g26775 (n14193, \a[25] , \a[57] );
  and g26776 (n14194, n7119, n14193);
  not g26777 (n_12841, n14192);
  not g26778 (n_12842, n14194);
  and g26779 (n14195, n_12841, n_12842);
  not g26780 (n_12843, n14191);
  not g26781 (n_12844, n14195);
  and g26782 (n14196, n_12843, n_12844);
  not g26783 (n_12845, n14196);
  and g26784 (n14197, n7119, n_12845);
  and g26785 (n14198, \a[27] , \a[55] );
  not g26786 (n_12846, n14193);
  not g26787 (n_12847, n14198);
  and g26788 (n14199, n_12846, n_12847);
  and g26789 (n14200, n_12843, n_12845);
  not g26790 (n_12848, n14199);
  and g26791 (n14201, n_12848, n14200);
  not g26792 (n_12849, n14197);
  not g26793 (n_12850, n14201);
  and g26794 (n14202, n_12849, n_12850);
  not g26795 (n_12851, n14190);
  not g26796 (n_12852, n14202);
  and g26797 (n14203, n_12851, n_12852);
  not g26798 (n_12853, n14203);
  and g26799 (n14204, n_12851, n_12853);
  and g26800 (n14205, n_12852, n_12853);
  not g26801 (n_12854, n14204);
  not g26802 (n_12855, n14205);
  and g26803 (n14206, n_12854, n_12855);
  and g26804 (n14207, n_12711, n_12715);
  and g26805 (n14208, n14206, n14207);
  not g26806 (n_12856, n14206);
  not g26807 (n_12857, n14207);
  and g26808 (n14209, n_12856, n_12857);
  not g26809 (n_12858, n14208);
  not g26810 (n_12859, n14209);
  and g26811 (n14210, n_12858, n_12859);
  and g26812 (n14211, n_12699, n14034);
  not g26813 (n_12860, n14211);
  and g26814 (n14212, n_12697, n_12860);
  and g26815 (n14213, n_12719, n_12722);
  not g26816 (n_12861, n14212);
  not g26817 (n_12862, n14213);
  and g26818 (n14214, n_12861, n_12862);
  not g26819 (n_12863, n14214);
  and g26820 (n14215, n_12861, n_12863);
  and g26821 (n14216, n_12862, n_12863);
  not g26822 (n_12864, n14215);
  not g26823 (n_12865, n14216);
  and g26824 (n14217, n_12864, n_12865);
  not g26825 (n_12866, n14217);
  and g26826 (n14218, n14210, n_12866);
  not g26827 (n_12867, n14210);
  and g26828 (n14219, n_12867, n14217);
  not g26829 (n_12868, n14189);
  not g26830 (n_12869, n14219);
  and g26831 (n14220, n_12868, n_12869);
  not g26832 (n_12870, n14218);
  and g26833 (n14221, n_12870, n14220);
  not g26834 (n_12871, n14221);
  and g26835 (n14222, n_12868, n_12871);
  and g26836 (n14223, n_12869, n_12871);
  and g26837 (n14224, n_12870, n14223);
  not g26838 (n_12872, n14222);
  not g26839 (n_12873, n14224);
  and g26840 (n14225, n_12872, n_12873);
  and g26841 (n14226, n_12580, n_12624);
  and g26842 (n14227, n13893, n14013);
  not g26843 (n_12874, n13893);
  not g26844 (n_12875, n14013);
  and g26845 (n14228, n_12874, n_12875);
  not g26846 (n_12876, n14227);
  not g26847 (n_12877, n14228);
  and g26848 (n14229, n_12876, n_12877);
  not g26849 (n_12878, n14229);
  and g26850 (n14230, n13945, n_12878);
  not g26851 (n_12879, n13945);
  and g26852 (n14231, n_12879, n14229);
  not g26853 (n_12880, n14230);
  not g26854 (n_12881, n14231);
  and g26855 (n14232, n_12880, n_12881);
  and g26856 (n14233, n13877, n13909);
  not g26857 (n_12882, n13877);
  not g26858 (n_12883, n13909);
  and g26859 (n14234, n_12882, n_12883);
  not g26860 (n_12884, n14233);
  not g26861 (n_12885, n14234);
  and g26862 (n14235, n_12884, n_12885);
  not g26863 (n_12886, n14235);
  and g26864 (n14236, n13927, n_12886);
  not g26865 (n_12887, n13927);
  and g26866 (n14237, n_12887, n14235);
  not g26867 (n_12888, n14236);
  not g26868 (n_12889, n14237);
  and g26869 (n14238, n_12888, n_12889);
  and g26870 (n14239, n_12603, n_12618);
  not g26871 (n_12890, n14238);
  and g26872 (n14240, n_12890, n14239);
  not g26873 (n_12891, n14239);
  and g26874 (n14241, n14238, n_12891);
  not g26875 (n_12892, n14240);
  not g26876 (n_12893, n14241);
  and g26877 (n14242, n_12892, n_12893);
  and g26878 (n14243, n14232, n14242);
  not g26879 (n_12894, n14232);
  not g26880 (n_12895, n14242);
  and g26881 (n14244, n_12894, n_12895);
  not g26882 (n_12896, n14243);
  not g26883 (n_12897, n14244);
  and g26884 (n14245, n_12896, n_12897);
  not g26885 (n_12898, n14245);
  and g26886 (n14246, n14226, n_12898);
  not g26887 (n_12899, n14226);
  and g26888 (n14247, n_12899, n14245);
  not g26889 (n_12900, n14246);
  not g26890 (n_12901, n14247);
  and g26891 (n14248, n_12900, n_12901);
  and g26892 (n14249, n_12671, n_12683);
  and g26893 (n14250, n_12562, n_12574);
  and g26894 (n14251, n14249, n14250);
  not g26895 (n_12902, n14249);
  not g26896 (n_12903, n14250);
  and g26897 (n14252, n_12902, n_12903);
  not g26898 (n_12904, n14251);
  not g26899 (n_12905, n14252);
  and g26900 (n14253, n_12904, n_12905);
  not g26901 (n_12906, n13863);
  and g26902 (n14254, n12547, n_12906);
  not g26903 (n_12907, n12547);
  and g26904 (n14255, n_12907, n13863);
  not g26905 (n_12908, n14254);
  not g26906 (n_12909, n14255);
  and g26907 (n14256, n_12908, n_12909);
  not g26908 (n_12910, n14256);
  and g26909 (n14257, n13977, n_12910);
  not g26910 (n_12911, n13977);
  and g26911 (n14258, n_12911, n14256);
  not g26912 (n_12912, n14257);
  not g26913 (n_12913, n14258);
  and g26914 (n14259, n_12912, n_12913);
  and g26915 (n14260, n14253, n14259);
  not g26916 (n_12914, n14253);
  not g26917 (n_12915, n14259);
  and g26918 (n14261, n_12914, n_12915);
  not g26919 (n_12916, n14260);
  not g26920 (n_12917, n14261);
  and g26921 (n14262, n_12916, n_12917);
  and g26922 (n14263, n14248, n14262);
  not g26923 (n_12918, n14248);
  not g26924 (n_12919, n14262);
  and g26925 (n14264, n_12918, n_12919);
  not g26926 (n_12920, n14263);
  not g26927 (n_12921, n14264);
  and g26928 (n14265, n_12920, n_12921);
  not g26929 (n_12922, n14225);
  not g26930 (n_12923, n14265);
  and g26931 (n14266, n_12922, n_12923);
  and g26932 (n14267, n14225, n14265);
  not g26933 (n_12924, n14266);
  not g26934 (n_12925, n14267);
  and g26935 (n14268, n_12924, n_12925);
  not g26936 (n_12926, n14188);
  not g26937 (n_12927, n14268);
  and g26938 (n14269, n_12926, n_12927);
  not g26939 (n_12928, n14269);
  and g26940 (n14270, n_12926, n_12928);
  and g26941 (n14271, n_12927, n_12928);
  not g26942 (n_12929, n14270);
  not g26943 (n_12930, n14271);
  and g26944 (n14272, n_12929, n_12930);
  not g26945 (n_12931, n14076);
  not g26946 (n_12932, n14272);
  and g26947 (n14273, n_12931, n_12932);
  and g26948 (n14274, n14076, n14272);
  not g26949 (n_12933, n14273);
  not g26950 (n_12934, n14274);
  and g26951 (n14275, n_12933, n_12934);
  not g26952 (n_12935, n14075);
  and g26953 (n14276, n_12935, n14275);
  not g26954 (n_12936, n14275);
  and g26955 (n14277, n14075, n_12936);
  not g26956 (n_12937, n14276);
  not g26957 (n_12938, n14277);
  and g26958 (\asquared[83] , n_12937, n_12938);
  and g26959 (n14279, n_12838, n_12928);
  and g26960 (n14280, n_12788, n_12826);
  and g26961 (n14281, n_12893, n_12896);
  not g26962 (n_12939, n14280);
  not g26963 (n_12940, n14281);
  and g26964 (n14282, n_12939, n_12940);
  not g26965 (n_12941, n14282);
  and g26966 (n14283, n_12939, n_12941);
  and g26967 (n14284, n_12940, n_12941);
  not g26968 (n_12942, n14283);
  not g26969 (n_12943, n14284);
  and g26970 (n14285, n_12942, n_12943);
  and g26971 (n14286, n14119, n14166);
  not g26972 (n_12944, n14119);
  not g26973 (n_12945, n14166);
  and g26974 (n14287, n_12944, n_12945);
  not g26975 (n_12946, n14286);
  not g26976 (n_12947, n14287);
  and g26977 (n14288, n_12946, n_12947);
  not g26978 (n_12948, n14288);
  and g26979 (n14289, n14139, n_12948);
  not g26980 (n_12949, n14139);
  and g26981 (n14290, n_12949, n14288);
  not g26982 (n_12950, n14289);
  not g26983 (n_12951, n14290);
  and g26984 (n14291, n_12950, n_12951);
  and g26985 (n14292, n14089, n14102);
  not g26986 (n_12952, n14089);
  not g26987 (n_12953, n14102);
  and g26988 (n14293, n_12952, n_12953);
  not g26989 (n_12954, n14292);
  not g26990 (n_12955, n14293);
  and g26991 (n14294, n_12954, n_12955);
  not g26992 (n_12956, n14294);
  and g26993 (n14295, n14200, n_12956);
  not g26994 (n_12957, n14200);
  and g26995 (n14296, n_12957, n14294);
  not g26996 (n_12958, n14295);
  not g26997 (n_12959, n14296);
  and g26998 (n14297, n_12958, n_12959);
  and g26999 (n14298, n_12805, n_12820);
  not g27000 (n_12960, n14297);
  and g27001 (n14299, n_12960, n14298);
  not g27002 (n_12961, n14298);
  and g27003 (n14300, n14297, n_12961);
  not g27004 (n_12962, n14299);
  not g27005 (n_12963, n14300);
  and g27006 (n14301, n_12962, n_12963);
  and g27007 (n14302, n14291, n14301);
  not g27008 (n_12964, n14291);
  not g27009 (n_12965, n14301);
  and g27010 (n14303, n_12964, n_12965);
  not g27011 (n_12966, n14302);
  not g27012 (n_12967, n14303);
  and g27013 (n14304, n_12966, n_12967);
  not g27014 (n_12968, n14285);
  and g27015 (n14305, n_12968, n14304);
  not g27016 (n_12969, n14305);
  and g27017 (n14306, n_12968, n_12969);
  and g27018 (n14307, n14304, n_12969);
  not g27019 (n_12970, n14306);
  not g27020 (n_12971, n14307);
  and g27021 (n14308, n_12970, n_12971);
  and g27022 (n14309, n_12828, n_12833);
  and g27023 (n14310, n_12877, n_12881);
  and g27024 (n14311, n_12885, n_12889);
  and g27025 (n14312, n14310, n14311);
  not g27026 (n_12972, n14310);
  not g27027 (n_12973, n14311);
  and g27028 (n14313, n_12972, n_12973);
  not g27029 (n_12974, n14312);
  not g27030 (n_12975, n14313);
  and g27031 (n14314, n_12974, n_12975);
  and g27032 (n14315, n_12767, n_12782);
  not g27033 (n_12976, n14314);
  and g27034 (n14316, n_12976, n14315);
  not g27035 (n_12977, n14315);
  and g27036 (n14317, n14314, n_12977);
  not g27037 (n_12978, n14316);
  not g27038 (n_12979, n14317);
  and g27039 (n14318, n_12978, n_12979);
  and g27040 (n14319, n1666, n9509);
  not g27041 (n_12980, n14319);
  and g27042 (n14320, \a[59] , n_12980);
  and g27043 (n14321, \a[24] , n14320);
  and g27044 (n14322, \a[60] , n_12980);
  and g27045 (n14323, \a[23] , n14322);
  not g27046 (n_12981, n14321);
  not g27047 (n_12982, n14323);
  and g27048 (n14324, n_12981, n_12982);
  not g27049 (n_12983, n14151);
  not g27050 (n_12984, n14324);
  and g27051 (n14325, n_12983, n_12984);
  not g27052 (n_12985, n14325);
  and g27053 (n14326, n_12983, n_12985);
  and g27054 (n14327, n_12984, n_12985);
  not g27055 (n_12986, n14326);
  not g27056 (n_12987, n14327);
  and g27057 (n14328, n_12986, n_12987);
  and g27058 (n14329, n3110, n7697);
  and g27059 (n14330, n2865, n7433);
  and g27060 (n14331, \a[31] , \a[55] );
  and g27061 (n14332, n13756, n14331);
  not g27062 (n_12988, n14330);
  not g27063 (n_12989, n14332);
  and g27064 (n14333, n_12988, n_12989);
  not g27065 (n_12990, n14329);
  not g27066 (n_12991, n14333);
  and g27067 (n14334, n_12990, n_12991);
  not g27068 (n_12992, n14334);
  and g27069 (n14335, \a[52] , n_12992);
  and g27070 (n14336, \a[31] , n14335);
  and g27071 (n14337, \a[28] , \a[55] );
  and g27072 (n14338, \a[30] , \a[53] );
  not g27073 (n_12993, n14337);
  not g27074 (n_12994, n14338);
  and g27075 (n14339, n_12993, n_12994);
  and g27076 (n14340, n_12990, n_12992);
  not g27077 (n_12995, n14339);
  and g27078 (n14341, n_12995, n14340);
  not g27079 (n_12996, n14336);
  not g27080 (n_12997, n14341);
  and g27081 (n14342, n_12996, n_12997);
  not g27082 (n_12998, n14328);
  not g27083 (n_12999, n14342);
  and g27084 (n14343, n_12998, n_12999);
  not g27085 (n_13000, n14343);
  and g27086 (n14344, n_12998, n_13000);
  and g27087 (n14345, n_12999, n_13000);
  not g27088 (n_13001, n14344);
  not g27089 (n_13002, n14345);
  and g27090 (n14346, n_13001, n_13002);
  and g27091 (n14347, n_12908, n_12913);
  and g27092 (n14348, n14346, n14347);
  not g27093 (n_13003, n14346);
  not g27094 (n_13004, n14347);
  and g27095 (n14349, n_13003, n_13004);
  not g27096 (n_13005, n14348);
  not g27097 (n_13006, n14349);
  and g27098 (n14350, n_13005, n_13006);
  and g27099 (n14351, n_12905, n_12916);
  not g27100 (n_13007, n14351);
  and g27101 (n14352, n14350, n_13007);
  not g27102 (n_13008, n14350);
  and g27103 (n14353, n_13008, n14351);
  not g27104 (n_13009, n14352);
  not g27105 (n_13010, n14353);
  and g27106 (n14354, n_13009, n_13010);
  and g27107 (n14355, n14318, n14354);
  not g27108 (n_13011, n14318);
  not g27109 (n_13012, n14354);
  and g27110 (n14356, n_13011, n_13012);
  not g27111 (n_13013, n14355);
  not g27112 (n_13014, n14356);
  and g27113 (n14357, n_13013, n_13014);
  not g27114 (n_13015, n14309);
  and g27115 (n14358, n_13015, n14357);
  not g27116 (n_13016, n14357);
  and g27117 (n14359, n14309, n_13016);
  not g27118 (n_13017, n14358);
  not g27119 (n_13018, n14359);
  and g27120 (n14360, n_13017, n_13018);
  and g27121 (n14361, n14308, n14360);
  not g27122 (n_13019, n14308);
  not g27123 (n_13020, n14360);
  and g27124 (n14362, n_13019, n_13020);
  not g27125 (n_13021, n14361);
  not g27126 (n_13022, n14362);
  and g27127 (n14363, n_13021, n_13022);
  and g27128 (n14364, n_12922, n14265);
  not g27129 (n_13023, n14364);
  and g27130 (n14365, n_12871, n_13023);
  and g27131 (n14366, n_12901, n_12920);
  and g27132 (n14367, n_12863, n_12870);
  and g27133 (n14368, \a[42] , \a[62] );
  and g27134 (n14369, \a[21] , n14368);
  not g27135 (n_13024, n14369);
  and g27136 (n14370, n5344, n_13024);
  not g27137 (n_13025, n14370);
  and g27138 (n14371, n_13024, n_13025);
  and g27139 (n14372, \a[21] , \a[62] );
  not g27140 (n_13026, \a[42] );
  not g27141 (n_13027, n14372);
  and g27142 (n14373, n_13026, n_13027);
  not g27143 (n_13028, n14373);
  and g27144 (n14374, n14371, n_13028);
  and g27145 (n14375, n5344, n_13025);
  not g27146 (n_13029, n14374);
  not g27147 (n_13030, n14375);
  and g27148 (n14376, n_13029, n_13030);
  and g27149 (n14377, \a[39] , \a[44] );
  and g27150 (n14378, \a[40] , \a[43] );
  not g27151 (n_13031, n14377);
  not g27152 (n_13032, n14378);
  and g27153 (n14379, n_13031, n_13032);
  and g27154 (n14380, n4171, n5296);
  not g27155 (n_13033, n14380);
  not g27158 (n_13034, n14379);
  not g27160 (n_13035, n14383);
  and g27161 (n14384, \a[54] , n_13035);
  and g27162 (n14385, \a[29] , n14384);
  and g27163 (n14386, n_13033, n_13035);
  and g27164 (n14387, n_13034, n14386);
  not g27165 (n_13036, n14385);
  not g27166 (n_13037, n14387);
  and g27167 (n14388, n_13036, n_13037);
  not g27168 (n_13038, n14376);
  not g27169 (n_13039, n14388);
  and g27170 (n14389, n_13038, n_13039);
  not g27171 (n_13040, n14389);
  and g27172 (n14390, n_13038, n_13040);
  and g27173 (n14391, n_13039, n_13040);
  not g27174 (n_13041, n14390);
  not g27175 (n_13042, n14391);
  and g27176 (n14392, n_13041, n_13042);
  and g27177 (n14393, n3319, n6256);
  and g27178 (n14394, n2972, n5888);
  and g27179 (n14395, n4150, n6325);
  not g27180 (n_13043, n14394);
  not g27181 (n_13044, n14395);
  and g27182 (n14396, n_13043, n_13044);
  not g27183 (n_13045, n14393);
  not g27184 (n_13046, n14396);
  and g27185 (n14397, n_13045, n_13046);
  not g27186 (n_13047, n14397);
  and g27187 (n14398, \a[50] , n_13047);
  and g27188 (n14399, \a[33] , n14398);
  and g27189 (n14400, n_13045, n_13047);
  and g27190 (n14401, \a[34] , \a[49] );
  and g27191 (n14402, \a[35] , \a[48] );
  not g27192 (n_13048, n14401);
  not g27193 (n_13049, n14402);
  and g27194 (n14403, n_13048, n_13049);
  not g27195 (n_13050, n14403);
  and g27196 (n14404, n14400, n_13050);
  not g27197 (n_13051, n14399);
  not g27198 (n_13052, n14404);
  and g27199 (n14405, n_13051, n_13052);
  not g27200 (n_13053, n14392);
  not g27201 (n_13054, n14405);
  and g27202 (n14406, n_13053, n_13054);
  not g27203 (n_13055, n14406);
  and g27204 (n14407, n_13053, n_13055);
  and g27205 (n14408, n_13054, n_13055);
  not g27206 (n_13056, n14407);
  not g27207 (n_13057, n14408);
  and g27208 (n14409, n_13056, n_13057);
  and g27209 (n14410, n_12853, n_12859);
  and g27210 (n14411, n14409, n14410);
  not g27211 (n_13058, n14409);
  not g27212 (n_13059, n14410);
  and g27213 (n14412, n_13058, n_13059);
  not g27214 (n_13060, n14411);
  not g27215 (n_13061, n14412);
  and g27216 (n14413, n_13060, n_13061);
  and g27217 (n14414, \a[26] , \a[57] );
  and g27218 (n14415, \a[32] , \a[51] );
  not g27219 (n_13062, n14414);
  not g27220 (n_13063, n14415);
  and g27221 (n14416, n_13062, n_13063);
  and g27222 (n14417, \a[51] , \a[57] );
  and g27223 (n14418, n3266, n14417);
  and g27224 (n14419, n2463, n8436);
  and g27225 (n14420, \a[32] , \a[58] );
  and g27226 (n14421, n12844, n14420);
  not g27227 (n_13064, n14419);
  not g27228 (n_13065, n14421);
  and g27229 (n14422, n_13064, n_13065);
  not g27230 (n_13066, n14418);
  not g27231 (n_13067, n14422);
  and g27232 (n14423, n_13066, n_13067);
  not g27233 (n_13068, n14423);
  and g27234 (n14424, n_13066, n_13068);
  not g27235 (n_13069, n14416);
  and g27236 (n14425, n_13069, n14424);
  and g27237 (n14426, \a[58] , n_13068);
  and g27238 (n14427, \a[25] , n14426);
  not g27239 (n_13070, n14425);
  not g27240 (n_13071, n14427);
  and g27241 (n14428, n_13070, n_13071);
  and g27242 (n14429, n4565, n5560);
  and g27243 (n14430, n3530, n5250);
  and g27244 (n14431, n3687, n5666);
  not g27245 (n_13072, n14430);
  not g27246 (n_13073, n14431);
  and g27247 (n14432, n_13072, n_13073);
  not g27248 (n_13074, n14429);
  not g27249 (n_13075, n14432);
  and g27250 (n14433, n_13074, n_13075);
  not g27251 (n_13076, n14433);
  and g27252 (n14434, \a[47] , n_13076);
  and g27253 (n14435, \a[36] , n14434);
  and g27254 (n14436, n_13074, n_13076);
  and g27255 (n14437, \a[37] , \a[46] );
  and g27256 (n14438, \a[38] , \a[45] );
  not g27257 (n_13077, n14437);
  not g27258 (n_13078, n14438);
  and g27259 (n14439, n_13077, n_13078);
  not g27260 (n_13079, n14439);
  and g27261 (n14440, n14436, n_13079);
  not g27262 (n_13080, n14435);
  not g27263 (n_13081, n14440);
  and g27264 (n14441, n_13080, n_13081);
  not g27265 (n_13082, n14428);
  not g27266 (n_13083, n14441);
  and g27267 (n14442, n_13082, n_13083);
  not g27268 (n_13084, n14442);
  and g27269 (n14443, n_13082, n_13084);
  and g27270 (n14444, n_13083, n_13084);
  not g27271 (n_13085, n14443);
  not g27272 (n_13086, n14444);
  and g27273 (n14445, n_13085, n_13086);
  and g27274 (n14446, \a[20] , \a[63] );
  and g27275 (n14447, \a[22] , \a[61] );
  not g27276 (n_13087, n14446);
  not g27277 (n_13088, n14447);
  and g27278 (n14448, n_13087, n_13088);
  and g27279 (n14449, n1693, n9909);
  not g27280 (n_13089, n14449);
  and g27281 (n14450, n13458, n_13089);
  not g27282 (n_13090, n14448);
  and g27283 (n14451, n_13090, n14450);
  not g27284 (n_13091, n14451);
  and g27285 (n14452, n13458, n_13091);
  and g27286 (n14453, n_13089, n_13091);
  and g27287 (n14454, n_13090, n14453);
  not g27288 (n_13092, n14452);
  not g27289 (n_13093, n14454);
  and g27290 (n14455, n_13092, n_13093);
  not g27291 (n_13094, n14445);
  not g27292 (n_13095, n14455);
  and g27293 (n14456, n_13094, n_13095);
  not g27294 (n_13096, n14456);
  and g27295 (n14457, n_13094, n_13096);
  and g27296 (n14458, n_13095, n_13096);
  not g27297 (n_13097, n14457);
  not g27298 (n_13098, n14458);
  and g27299 (n14459, n_13097, n_13098);
  not g27300 (n_13099, n14413);
  and g27301 (n14460, n_13099, n14459);
  not g27302 (n_13100, n14459);
  and g27303 (n14461, n14413, n_13100);
  not g27304 (n_13101, n14460);
  not g27305 (n_13102, n14461);
  and g27306 (n14462, n_13101, n_13102);
  not g27307 (n_13103, n14367);
  and g27308 (n14463, n_13103, n14462);
  not g27309 (n_13104, n14462);
  and g27310 (n14464, n14367, n_13104);
  not g27311 (n_13105, n14463);
  not g27312 (n_13106, n14464);
  and g27313 (n14465, n_13105, n_13106);
  not g27314 (n_13107, n14366);
  and g27315 (n14466, n_13107, n14465);
  not g27316 (n_13108, n14465);
  and g27317 (n14467, n14366, n_13108);
  not g27318 (n_13109, n14466);
  not g27319 (n_13110, n14467);
  and g27320 (n14468, n_13109, n_13110);
  not g27321 (n_13111, n14365);
  and g27322 (n14469, n_13111, n14468);
  not g27323 (n_13112, n14468);
  and g27324 (n14470, n14365, n_13112);
  not g27325 (n_13113, n14469);
  not g27326 (n_13114, n14470);
  and g27327 (n14471, n_13113, n_13114);
  not g27328 (n_13115, n14363);
  and g27329 (n14472, n_13115, n14471);
  not g27330 (n_13116, n14472);
  and g27331 (n14473, n14471, n_13116);
  and g27332 (n14474, n_13115, n_13116);
  not g27333 (n_13117, n14473);
  not g27334 (n_13118, n14474);
  and g27335 (n14475, n_13117, n_13118);
  not g27336 (n_13119, n14279);
  not g27337 (n_13120, n14475);
  and g27338 (n14476, n_13119, n_13120);
  and g27339 (n14477, n14279, n14475);
  not g27340 (n_13121, n14476);
  not g27341 (n_13122, n14477);
  and g27342 (n14478, n_13121, n_13122);
  and g27343 (n14479, n_12935, n_12934);
  not g27344 (n_13123, n14479);
  and g27345 (n14480, n_12933, n_13123);
  not g27346 (n_13124, n14478);
  and g27347 (n14481, n_13124, n14480);
  not g27348 (n_13125, n14480);
  and g27349 (n14482, n14478, n_13125);
  not g27350 (n_13126, n14481);
  not g27351 (n_13127, n14482);
  and g27352 (\asquared[84] , n_13126, n_13127);
  and g27353 (n14484, n_13122, n_13125);
  not g27354 (n_13128, n14484);
  and g27355 (n14485, n_13121, n_13128);
  and g27356 (n14486, n_13113, n_13116);
  and g27357 (n14487, n_13019, n14360);
  not g27358 (n_13129, n14487);
  and g27359 (n14488, n_13017, n_13129);
  and g27360 (n14489, n_12980, n_12985);
  and g27361 (n14490, n14453, n14489);
  not g27362 (n_13130, n14453);
  not g27363 (n_13131, n14489);
  and g27364 (n14491, n_13130, n_13131);
  not g27365 (n_13132, n14490);
  not g27366 (n_13133, n14491);
  and g27367 (n14492, n_13132, n_13133);
  and g27368 (n14493, \a[31] , \a[53] );
  and g27369 (n14494, \a[32] , \a[52] );
  not g27370 (n_13134, n14493);
  not g27371 (n_13135, n14494);
  and g27372 (n14495, n_13134, n_13135);
  and g27373 (n14496, n3812, n7433);
  not g27374 (n_13136, n14496);
  and g27375 (n14497, n12603, n_13136);
  not g27376 (n_13137, n14495);
  and g27377 (n14498, n_13137, n14497);
  not g27378 (n_13138, n14498);
  and g27379 (n14499, n12603, n_13138);
  and g27380 (n14500, n_13136, n_13138);
  and g27381 (n14501, n_13137, n14500);
  not g27382 (n_13139, n14499);
  not g27383 (n_13140, n14501);
  and g27384 (n14502, n_13139, n_13140);
  not g27385 (n_13141, n14502);
  and g27386 (n14503, n14492, n_13141);
  not g27387 (n_13142, n14503);
  and g27388 (n14504, n14492, n_13142);
  and g27389 (n14505, n_13141, n_13142);
  not g27390 (n_13143, n14504);
  not g27391 (n_13144, n14505);
  and g27392 (n14506, n_13143, n_13144);
  and g27393 (n14507, n_13000, n_13006);
  and g27394 (n14508, n14506, n14507);
  not g27395 (n_13145, n14506);
  not g27396 (n_13146, n14507);
  and g27397 (n14509, n_13145, n_13146);
  not g27398 (n_13147, n14508);
  not g27399 (n_13148, n14509);
  and g27400 (n14510, n_13147, n_13148);
  and g27401 (n14511, n_12975, n_12979);
  not g27402 (n_13149, n14510);
  and g27403 (n14512, n_13149, n14511);
  not g27404 (n_13150, n14511);
  and g27405 (n14513, n14510, n_13150);
  not g27406 (n_13151, n14512);
  not g27407 (n_13152, n14513);
  and g27408 (n14514, n_13151, n_13152);
  and g27409 (n14515, n_13009, n_13013);
  not g27410 (n_13153, n14514);
  and g27411 (n14516, n_13153, n14515);
  not g27412 (n_13154, n14515);
  and g27413 (n14517, n14514, n_13154);
  not g27414 (n_13155, n14516);
  not g27415 (n_13156, n14517);
  and g27416 (n14518, n_13155, n_13156);
  and g27417 (n14519, n1919, n9721);
  and g27418 (n14520, n1367, n9909);
  and g27419 (n14521, n1574, n9792);
  not g27420 (n_13157, n14520);
  not g27421 (n_13158, n14521);
  and g27422 (n14522, n_13157, n_13158);
  not g27423 (n_13159, n14519);
  not g27424 (n_13160, n14522);
  and g27425 (n14523, n_13159, n_13160);
  not g27426 (n_13161, n14523);
  and g27427 (n14524, n_13159, n_13161);
  and g27428 (n14525, \a[22] , \a[62] );
  and g27429 (n14526, \a[23] , \a[61] );
  not g27430 (n_13162, n14525);
  not g27431 (n_13163, n14526);
  and g27432 (n14527, n_13162, n_13163);
  not g27433 (n_13164, n14527);
  and g27434 (n14528, n14524, n_13164);
  and g27435 (n14529, \a[63] , n_13161);
  and g27436 (n14530, \a[21] , n14529);
  not g27437 (n_13165, n14528);
  not g27438 (n_13166, n14530);
  and g27439 (n14531, n_13165, n_13166);
  and g27440 (n14532, \a[24] , \a[60] );
  and g27441 (n14533, \a[25] , \a[59] );
  not g27442 (n_13167, n14532);
  not g27443 (n_13168, n14533);
  and g27444 (n14534, n_13167, n_13168);
  and g27445 (n14535, n1904, n9509);
  not g27446 (n_13169, n14535);
  not g27449 (n_13170, n14534);
  not g27451 (n_13171, n14538);
  and g27452 (n14539, \a[51] , n_13171);
  and g27453 (n14540, \a[33] , n14539);
  and g27454 (n14541, n_13169, n_13171);
  and g27455 (n14542, n_13170, n14541);
  not g27456 (n_13172, n14540);
  not g27457 (n_13173, n14542);
  and g27458 (n14543, n_13172, n_13173);
  not g27459 (n_13174, n14531);
  not g27460 (n_13175, n14543);
  and g27461 (n14544, n_13174, n_13175);
  not g27462 (n_13176, n14544);
  and g27463 (n14545, n_13174, n_13176);
  and g27464 (n14546, n_13175, n_13176);
  not g27465 (n_13177, n14545);
  not g27466 (n_13178, n14546);
  and g27467 (n14547, n_13177, n_13178);
  and g27468 (n14548, n3828, n6256);
  and g27469 (n14549, n4595, n5888);
  and g27470 (n14550, n3319, n6325);
  not g27471 (n_13179, n14549);
  not g27472 (n_13180, n14550);
  and g27473 (n14551, n_13179, n_13180);
  not g27474 (n_13181, n14548);
  not g27475 (n_13182, n14551);
  and g27476 (n14552, n_13181, n_13182);
  not g27477 (n_13183, n14552);
  and g27478 (n14553, \a[50] , n_13183);
  and g27479 (n14554, \a[34] , n14553);
  and g27480 (n14555, n_13181, n_13183);
  and g27481 (n14556, \a[35] , \a[49] );
  and g27482 (n14557, \a[36] , \a[48] );
  not g27483 (n_13184, n14556);
  not g27484 (n_13185, n14557);
  and g27485 (n14558, n_13184, n_13185);
  not g27486 (n_13186, n14558);
  and g27487 (n14559, n14555, n_13186);
  not g27488 (n_13187, n14554);
  not g27489 (n_13188, n14559);
  and g27490 (n14560, n_13187, n_13188);
  not g27491 (n_13189, n14547);
  not g27492 (n_13190, n14560);
  and g27493 (n14561, n_13189, n_13190);
  not g27494 (n_13191, n14561);
  and g27495 (n14562, n_13189, n_13191);
  and g27496 (n14563, n_13190, n_13191);
  not g27497 (n_13192, n14562);
  not g27498 (n_13193, n14563);
  and g27499 (n14564, n_13192, n_13193);
  and g27500 (n14565, \a[29] , \a[55] );
  and g27501 (n14566, \a[38] , \a[46] );
  not g27502 (n_13194, n14565);
  not g27503 (n_13195, n14566);
  and g27504 (n14567, n_13194, n_13195);
  and g27505 (n14568, n2334, n9161);
  and g27506 (n14569, \a[38] , \a[56] );
  and g27507 (n14570, n12377, n14569);
  not g27508 (n_13196, n14568);
  not g27509 (n_13197, n14570);
  and g27510 (n14571, n_13196, n_13197);
  and g27511 (n14572, n14565, n14566);
  not g27512 (n_13198, n14571);
  not g27513 (n_13199, n14572);
  and g27514 (n14573, n_13198, n_13199);
  not g27515 (n_13200, n14573);
  and g27516 (n14574, n_13199, n_13200);
  not g27517 (n_13201, n14567);
  and g27518 (n14575, n_13201, n14574);
  and g27519 (n14576, \a[56] , n_13200);
  and g27520 (n14577, \a[28] , n14576);
  not g27521 (n_13202, n14575);
  not g27522 (n_13203, n14577);
  and g27523 (n14578, n_13202, n_13203);
  and g27524 (n14579, n5296, n5413);
  and g27525 (n14580, n3984, n4811);
  and g27526 (n14581, n4171, n5713);
  not g27527 (n_13204, n14580);
  not g27528 (n_13205, n14581);
  and g27529 (n14582, n_13204, n_13205);
  not g27530 (n_13206, n14579);
  not g27531 (n_13207, n14582);
  and g27532 (n14583, n_13206, n_13207);
  not g27533 (n_13208, n14583);
  and g27534 (n14584, \a[45] , n_13208);
  and g27535 (n14585, \a[39] , n14584);
  and g27536 (n14586, n_13206, n_13208);
  and g27537 (n14587, \a[40] , \a[44] );
  not g27538 (n_13209, n4807);
  not g27539 (n_13210, n14587);
  and g27540 (n14588, n_13209, n_13210);
  not g27541 (n_13211, n14588);
  and g27542 (n14589, n14586, n_13211);
  not g27543 (n_13212, n14585);
  not g27544 (n_13213, n14589);
  and g27545 (n14590, n_13212, n_13213);
  not g27546 (n_13214, n14578);
  not g27547 (n_13215, n14590);
  and g27548 (n14591, n_13214, n_13215);
  not g27549 (n_13216, n14591);
  and g27550 (n14592, n_13214, n_13216);
  and g27551 (n14593, n_13215, n_13216);
  not g27552 (n_13217, n14592);
  not g27553 (n_13218, n14593);
  and g27554 (n14594, n_13217, n_13218);
  and g27555 (n14595, \a[27] , \a[57] );
  and g27556 (n14596, \a[30] , \a[54] );
  not g27557 (n_13219, n14595);
  not g27558 (n_13220, n14596);
  and g27559 (n14597, n_13219, n_13220);
  and g27560 (n14598, \a[30] , \a[57] );
  and g27561 (n14599, n13969, n14598);
  not g27562 (n_13221, n14599);
  and g27563 (n14600, n14159, n_13221);
  not g27564 (n_13222, n14597);
  and g27565 (n14601, n_13222, n14600);
  not g27566 (n_13223, n14601);
  and g27567 (n14602, n14159, n_13223);
  and g27568 (n14603, n_13221, n_13223);
  and g27569 (n14604, n_13222, n14603);
  not g27570 (n_13224, n14602);
  not g27571 (n_13225, n14604);
  and g27572 (n14605, n_13224, n_13225);
  not g27573 (n_13226, n14594);
  not g27574 (n_13227, n14605);
  and g27575 (n14606, n_13226, n_13227);
  not g27576 (n_13228, n14606);
  and g27577 (n14607, n_13226, n_13228);
  and g27578 (n14608, n_13227, n_13228);
  not g27579 (n_13229, n14607);
  not g27580 (n_13230, n14608);
  and g27581 (n14609, n_13229, n_13230);
  not g27582 (n_13231, n14564);
  and g27583 (n14610, n_13231, n14609);
  not g27584 (n_13232, n14609);
  and g27585 (n14611, n14564, n_13232);
  not g27586 (n_13233, n14610);
  not g27587 (n_13234, n14611);
  and g27588 (n14612, n_13233, n_13234);
  and g27589 (n14613, n14400, n14436);
  not g27590 (n_13235, n14400);
  not g27591 (n_13236, n14436);
  and g27592 (n14614, n_13235, n_13236);
  not g27593 (n_13237, n14613);
  not g27594 (n_13238, n14614);
  and g27595 (n14615, n_13237, n_13238);
  not g27596 (n_13239, n14615);
  and g27597 (n14616, n14424, n_13239);
  not g27598 (n_13240, n14424);
  and g27599 (n14617, n_13240, n14615);
  not g27600 (n_13241, n14616);
  not g27601 (n_13242, n14617);
  and g27602 (n14618, n_13241, n_13242);
  and g27603 (n14619, n_12947, n_12951);
  and g27604 (n14620, n_12955, n_12959);
  and g27605 (n14621, n14619, n14620);
  not g27606 (n_13243, n14619);
  not g27607 (n_13244, n14620);
  and g27608 (n14622, n_13243, n_13244);
  not g27609 (n_13245, n14621);
  not g27610 (n_13246, n14622);
  and g27611 (n14623, n_13245, n_13246);
  and g27612 (n14624, n14618, n14623);
  not g27613 (n_13247, n14618);
  not g27614 (n_13248, n14623);
  and g27615 (n14625, n_13247, n_13248);
  not g27616 (n_13249, n14624);
  not g27617 (n_13250, n14625);
  and g27618 (n14626, n_13249, n_13250);
  not g27619 (n_13251, n14612);
  and g27620 (n14627, n_13251, n14626);
  not g27621 (n_13252, n14627);
  and g27622 (n14628, n_13251, n_13252);
  and g27623 (n14629, n14626, n_13252);
  not g27624 (n_13253, n14628);
  not g27625 (n_13254, n14629);
  and g27626 (n14630, n_13253, n_13254);
  not g27627 (n_13255, n14630);
  and g27628 (n14631, n14518, n_13255);
  not g27629 (n_13256, n14518);
  and g27630 (n14632, n_13256, n14630);
  not g27631 (n_13257, n14488);
  not g27632 (n_13258, n14632);
  and g27633 (n14633, n_13257, n_13258);
  not g27634 (n_13259, n14631);
  and g27635 (n14634, n_13259, n14633);
  not g27636 (n_13260, n14634);
  and g27637 (n14635, n_13257, n_13260);
  and g27638 (n14636, n_13258, n_13260);
  and g27639 (n14637, n_13259, n14636);
  not g27640 (n_13261, n14635);
  not g27641 (n_13262, n14637);
  and g27642 (n14638, n_13261, n_13262);
  and g27643 (n14639, n_13105, n_13109);
  and g27644 (n14640, n_12941, n_12969);
  and g27645 (n14641, n14639, n14640);
  not g27646 (n_13263, n14639);
  not g27647 (n_13264, n14640);
  and g27648 (n14642, n_13263, n_13264);
  not g27649 (n_13265, n14641);
  not g27650 (n_13266, n14642);
  and g27651 (n14643, n_13265, n_13266);
  and g27652 (n14644, n_13061, n_13102);
  and g27653 (n14645, n_12963, n_12966);
  not g27654 (n_13267, n14644);
  not g27655 (n_13268, n14645);
  and g27656 (n14646, n_13267, n_13268);
  not g27657 (n_13269, n14646);
  and g27658 (n14647, n_13267, n_13269);
  and g27659 (n14648, n_13268, n_13269);
  not g27660 (n_13270, n14647);
  not g27661 (n_13271, n14648);
  and g27662 (n14649, n_13270, n_13271);
  and g27663 (n14650, n14371, n14386);
  not g27664 (n_13272, n14371);
  not g27665 (n_13273, n14386);
  and g27666 (n14651, n_13272, n_13273);
  not g27667 (n_13274, n14650);
  not g27668 (n_13275, n14651);
  and g27669 (n14652, n_13274, n_13275);
  not g27670 (n_13276, n14652);
  and g27671 (n14653, n14340, n_13276);
  not g27672 (n_13277, n14340);
  and g27673 (n14654, n_13277, n14652);
  not g27674 (n_13278, n14653);
  not g27675 (n_13279, n14654);
  and g27676 (n14655, n_13278, n_13279);
  and g27677 (n14656, n_13084, n_13096);
  and g27678 (n14657, n_13040, n_13055);
  and g27679 (n14658, n14656, n14657);
  not g27680 (n_13280, n14656);
  not g27681 (n_13281, n14657);
  and g27682 (n14659, n_13280, n_13281);
  not g27683 (n_13282, n14658);
  not g27684 (n_13283, n14659);
  and g27685 (n14660, n_13282, n_13283);
  and g27686 (n14661, n14655, n14660);
  not g27687 (n_13284, n14655);
  not g27688 (n_13285, n14660);
  and g27689 (n14662, n_13284, n_13285);
  not g27690 (n_13286, n14661);
  not g27691 (n_13287, n14662);
  and g27692 (n14663, n_13286, n_13287);
  not g27693 (n_13288, n14649);
  and g27694 (n14664, n_13288, n14663);
  not g27695 (n_13289, n14664);
  and g27696 (n14665, n_13288, n_13289);
  and g27697 (n14666, n14663, n_13289);
  not g27698 (n_13290, n14665);
  not g27699 (n_13291, n14666);
  and g27700 (n14667, n_13290, n_13291);
  not g27701 (n_13292, n14667);
  and g27702 (n14668, n14643, n_13292);
  not g27703 (n_13293, n14643);
  and g27704 (n14669, n_13293, n14667);
  not g27705 (n_13294, n14638);
  not g27706 (n_13295, n14669);
  and g27707 (n14670, n_13294, n_13295);
  not g27708 (n_13296, n14668);
  and g27709 (n14671, n_13296, n14670);
  not g27710 (n_13297, n14671);
  and g27711 (n14672, n_13294, n_13297);
  and g27712 (n14673, n_13295, n_13297);
  and g27713 (n14674, n_13296, n14673);
  not g27714 (n_13298, n14672);
  not g27715 (n_13299, n14674);
  and g27716 (n14675, n_13298, n_13299);
  not g27717 (n_13300, n14486);
  not g27718 (n_13301, n14675);
  and g27719 (n14676, n_13300, n_13301);
  and g27720 (n14677, n14486, n14675);
  not g27721 (n_13302, n14676);
  not g27722 (n_13303, n14677);
  and g27723 (n14678, n_13302, n_13303);
  not g27724 (n_13304, n14485);
  and g27725 (n14679, n_13304, n14678);
  not g27726 (n_13305, n14678);
  and g27727 (n14680, n14485, n_13305);
  not g27728 (n_13306, n14679);
  not g27729 (n_13307, n14680);
  and g27730 (\asquared[85] , n_13306, n_13307);
  and g27731 (n14682, n_13304, n_13303);
  not g27732 (n_13308, n14682);
  and g27733 (n14683, n_13302, n_13308);
  and g27734 (n14684, n_13260, n_13297);
  and g27735 (n14685, n_13266, n_13296);
  and g27736 (n14686, \a[22] , \a[63] );
  and g27737 (n14687, \a[28] , \a[57] );
  not g27738 (n_13309, n14686);
  not g27739 (n_13310, n14687);
  and g27740 (n14688, n_13309, n_13310);
  and g27741 (n14689, n14686, n14687);
  not g27742 (n_13311, n14689);
  not g27745 (n_13312, n14688);
  not g27747 (n_13313, n14692);
  and g27748 (n14693, n_13311, n_13313);
  and g27749 (n14694, n_13312, n14693);
  and g27750 (n14695, \a[50] , n_13313);
  and g27751 (n14696, \a[35] , n14695);
  not g27752 (n_13314, n14694);
  not g27753 (n_13315, n14696);
  and g27754 (n14697, n_13314, n_13315);
  and g27755 (n14698, n4150, n6968);
  and g27756 (n14699, n4090, n7232);
  and g27757 (n14700, n3143, n7433);
  not g27758 (n_13316, n14699);
  not g27759 (n_13317, n14700);
  and g27760 (n14701, n_13316, n_13317);
  not g27761 (n_13318, n14698);
  not g27762 (n_13319, n14701);
  and g27763 (n14702, n_13318, n_13319);
  not g27764 (n_13320, n14702);
  and g27765 (n14703, \a[53] , n_13320);
  and g27766 (n14704, \a[32] , n14703);
  and g27767 (n14705, n_13318, n_13320);
  and g27768 (n14706, \a[33] , \a[52] );
  and g27769 (n14707, \a[34] , \a[51] );
  not g27770 (n_13321, n14706);
  not g27771 (n_13322, n14707);
  and g27772 (n14708, n_13321, n_13322);
  not g27773 (n_13323, n14708);
  and g27774 (n14709, n14705, n_13323);
  not g27775 (n_13324, n14704);
  not g27776 (n_13325, n14709);
  and g27777 (n14710, n_13324, n_13325);
  not g27778 (n_13326, n14697);
  not g27779 (n_13327, n14710);
  and g27780 (n14711, n_13326, n_13327);
  not g27781 (n_13328, n14711);
  and g27782 (n14712, n_13326, n_13328);
  and g27783 (n14713, n_13327, n_13328);
  not g27784 (n_13329, n14712);
  not g27785 (n_13330, n14713);
  and g27786 (n14714, n_13329, n_13330);
  and g27787 (n14715, n5413, n5713);
  and g27788 (n14716, n3984, n7747);
  and g27789 (n14717, n4171, n5560);
  not g27790 (n_13331, n14716);
  not g27791 (n_13332, n14717);
  and g27792 (n14718, n_13331, n_13332);
  not g27793 (n_13333, n14715);
  not g27794 (n_13334, n14718);
  and g27795 (n14719, n_13333, n_13334);
  not g27796 (n_13335, n14719);
  and g27797 (n14720, \a[46] , n_13335);
  and g27798 (n14721, \a[39] , n14720);
  and g27799 (n14722, n_13333, n_13335);
  and g27800 (n14723, \a[40] , \a[45] );
  and g27801 (n14724, \a[41] , \a[44] );
  not g27802 (n_13336, n14723);
  not g27803 (n_13337, n14724);
  and g27804 (n14725, n_13336, n_13337);
  not g27805 (n_13338, n14725);
  and g27806 (n14726, n14722, n_13338);
  not g27807 (n_13339, n14721);
  not g27808 (n_13340, n14726);
  and g27809 (n14727, n_13339, n_13340);
  not g27810 (n_13341, n14714);
  not g27811 (n_13342, n14727);
  and g27812 (n14728, n_13341, n_13342);
  not g27813 (n_13343, n14728);
  and g27814 (n14729, n_13341, n_13343);
  and g27815 (n14730, n_13342, n_13343);
  not g27816 (n_13344, n14729);
  not g27817 (n_13345, n14730);
  and g27818 (n14731, n_13344, n_13345);
  and g27819 (n14732, \a[43] , \a[62] );
  and g27820 (n14733, \a[23] , n14732);
  not g27821 (n_13346, n14733);
  and g27822 (n14734, n5018, n_13346);
  not g27823 (n_13347, n14734);
  and g27824 (n14735, n_13346, n_13347);
  and g27825 (n14736, \a[23] , \a[62] );
  not g27826 (n_13348, \a[43] );
  not g27827 (n_13349, n14736);
  and g27828 (n14737, n_13348, n_13349);
  not g27829 (n_13350, n14737);
  and g27830 (n14738, n14735, n_13350);
  and g27831 (n14739, n5018, n_13347);
  not g27832 (n_13351, n14738);
  not g27833 (n_13352, n14739);
  and g27834 (n14740, n_13351, n_13352);
  and g27835 (n14741, n4565, n6252);
  and g27836 (n14742, n3530, n6254);
  and g27837 (n14743, n3687, n6256);
  not g27838 (n_13353, n14742);
  not g27839 (n_13354, n14743);
  and g27840 (n14744, n_13353, n_13354);
  not g27841 (n_13355, n14741);
  not g27842 (n_13356, n14744);
  and g27843 (n14745, n_13355, n_13356);
  not g27844 (n_13357, n14745);
  and g27845 (n14746, \a[49] , n_13357);
  and g27846 (n14747, \a[36] , n14746);
  and g27847 (n14748, \a[37] , \a[48] );
  and g27848 (n14749, \a[38] , \a[47] );
  not g27849 (n_13358, n14748);
  not g27850 (n_13359, n14749);
  and g27851 (n14750, n_13358, n_13359);
  and g27852 (n14751, n_13355, n_13357);
  not g27853 (n_13360, n14750);
  and g27854 (n14752, n_13360, n14751);
  not g27855 (n_13361, n14747);
  not g27856 (n_13362, n14752);
  and g27857 (n14753, n_13361, n_13362);
  not g27858 (n_13363, n14740);
  not g27859 (n_13364, n14753);
  and g27860 (n14754, n_13363, n_13364);
  not g27861 (n_13365, n14754);
  and g27862 (n14755, n_13363, n_13365);
  and g27863 (n14756, n_13364, n_13365);
  not g27864 (n_13366, n14755);
  not g27865 (n_13367, n14756);
  and g27866 (n14757, n_13366, n_13367);
  and g27867 (n14758, n2865, n7701);
  and g27868 (n14759, n3452, n7421);
  and g27869 (n14760, n2617, n9161);
  not g27870 (n_13368, n14759);
  not g27871 (n_13369, n14760);
  and g27872 (n14761, n_13368, n_13369);
  not g27873 (n_13370, n14758);
  not g27874 (n_13371, n14761);
  and g27875 (n14762, n_13370, n_13371);
  not g27876 (n_13372, n14762);
  and g27877 (n14763, \a[56] , n_13372);
  and g27878 (n14764, \a[29] , n14763);
  and g27879 (n14765, n_13370, n_13372);
  and g27880 (n14766, \a[30] , \a[55] );
  and g27881 (n14767, \a[31] , \a[54] );
  not g27882 (n_13373, n14766);
  not g27883 (n_13374, n14767);
  and g27884 (n14768, n_13373, n_13374);
  not g27885 (n_13375, n14768);
  and g27886 (n14769, n14765, n_13375);
  not g27887 (n_13376, n14764);
  not g27888 (n_13377, n14769);
  and g27889 (n14770, n_13376, n_13377);
  not g27890 (n_13378, n14757);
  not g27891 (n_13379, n14770);
  and g27892 (n14771, n_13378, n_13379);
  not g27893 (n_13380, n14771);
  and g27894 (n14772, n_13378, n_13380);
  and g27895 (n14773, n_13379, n_13380);
  not g27896 (n_13381, n14772);
  not g27897 (n_13382, n14773);
  and g27898 (n14774, n_13381, n_13382);
  not g27899 (n_13383, n14731);
  and g27900 (n14775, n_13383, n14774);
  not g27901 (n_13384, n14774);
  and g27902 (n14776, n14731, n_13384);
  not g27903 (n_13385, n14775);
  not g27904 (n_13386, n14776);
  and g27905 (n14777, n_13385, n_13386);
  and g27906 (n14778, n_13283, n_13286);
  and g27907 (n14779, n14777, n14778);
  not g27908 (n_13387, n14777);
  not g27909 (n_13388, n14778);
  and g27910 (n14780, n_13387, n_13388);
  not g27911 (n_13389, n14779);
  not g27912 (n_13390, n14780);
  and g27913 (n14781, n_13389, n_13390);
  and g27914 (n14782, n_13246, n_13249);
  and g27915 (n14783, \a[24] , \a[61] );
  not g27916 (n_13391, n14586);
  and g27917 (n14784, n_13391, n14783);
  not g27918 (n_13392, n14783);
  and g27919 (n14785, n14586, n_13392);
  not g27920 (n_13393, n14784);
  not g27921 (n_13394, n14785);
  and g27922 (n14786, n_13393, n_13394);
  not g27923 (n_13395, n14786);
  and g27924 (n14787, n14574, n_13395);
  not g27925 (n_13396, n14574);
  and g27926 (n14788, n_13396, n14786);
  not g27927 (n_13397, n14787);
  not g27928 (n_13398, n14788);
  and g27929 (n14789, n_13397, n_13398);
  and g27930 (n14790, n14500, n14603);
  not g27931 (n_13399, n14500);
  not g27932 (n_13400, n14603);
  and g27933 (n14791, n_13399, n_13400);
  not g27934 (n_13401, n14790);
  not g27935 (n_13402, n14791);
  and g27936 (n14792, n_13401, n_13402);
  and g27937 (n14793, n2227, n8987);
  and g27938 (n14794, n2633, n10089);
  and g27939 (n14795, n2463, n9509);
  not g27940 (n_13403, n14794);
  not g27941 (n_13404, n14795);
  and g27942 (n14796, n_13403, n_13404);
  not g27943 (n_13405, n14793);
  not g27944 (n_13406, n14796);
  and g27945 (n14797, n_13405, n_13406);
  not g27946 (n_13407, n14797);
  and g27947 (n14798, \a[60] , n_13407);
  and g27948 (n14799, \a[25] , n14798);
  and g27949 (n14800, n_13405, n_13407);
  and g27950 (n14801, \a[27] , \a[58] );
  not g27951 (n_13408, n8311);
  not g27952 (n_13409, n14801);
  and g27953 (n14802, n_13408, n_13409);
  not g27954 (n_13410, n14802);
  and g27955 (n14803, n14800, n_13410);
  not g27956 (n_13411, n14799);
  not g27957 (n_13412, n14803);
  and g27958 (n14804, n_13411, n_13412);
  not g27959 (n_13413, n14804);
  and g27960 (n14805, n14792, n_13413);
  not g27961 (n_13414, n14805);
  and g27962 (n14806, n14792, n_13414);
  and g27963 (n14807, n_13413, n_13414);
  not g27964 (n_13415, n14806);
  not g27965 (n_13416, n14807);
  and g27966 (n14808, n_13415, n_13416);
  not g27967 (n_13417, n14808);
  and g27968 (n14809, n14789, n_13417);
  not g27969 (n_13418, n14789);
  and g27970 (n14810, n_13418, n14808);
  not g27971 (n_13419, n14782);
  not g27972 (n_13420, n14810);
  and g27973 (n14811, n_13419, n_13420);
  not g27974 (n_13421, n14809);
  and g27975 (n14812, n_13421, n14811);
  not g27976 (n_13422, n14812);
  and g27977 (n14813, n_13419, n_13422);
  and g27978 (n14814, n_13421, n_13422);
  and g27979 (n14815, n_13420, n14814);
  not g27980 (n_13423, n14813);
  not g27981 (n_13424, n14815);
  and g27982 (n14816, n_13423, n_13424);
  and g27983 (n14817, n14524, n14555);
  not g27984 (n_13425, n14524);
  not g27985 (n_13426, n14555);
  and g27986 (n14818, n_13425, n_13426);
  not g27987 (n_13427, n14817);
  not g27988 (n_13428, n14818);
  and g27989 (n14819, n_13427, n_13428);
  not g27990 (n_13429, n14819);
  and g27991 (n14820, n14541, n_13429);
  not g27992 (n_13430, n14541);
  and g27993 (n14821, n_13430, n14819);
  not g27994 (n_13431, n14820);
  not g27995 (n_13432, n14821);
  and g27996 (n14822, n_13431, n_13432);
  and g27997 (n14823, n_13216, n_13228);
  and g27998 (n14824, n_13176, n_13191);
  and g27999 (n14825, n14823, n14824);
  not g28000 (n_13433, n14823);
  not g28001 (n_13434, n14824);
  and g28002 (n14826, n_13433, n_13434);
  not g28003 (n_13435, n14825);
  not g28004 (n_13436, n14826);
  and g28005 (n14827, n_13435, n_13436);
  and g28006 (n14828, n14822, n14827);
  not g28007 (n_13437, n14822);
  not g28008 (n_13438, n14827);
  and g28009 (n14829, n_13437, n_13438);
  not g28010 (n_13439, n14828);
  not g28011 (n_13440, n14829);
  and g28012 (n14830, n_13439, n_13440);
  not g28013 (n_13441, n14816);
  and g28014 (n14831, n_13441, n14830);
  not g28015 (n_13442, n14831);
  and g28016 (n14832, n_13441, n_13442);
  and g28017 (n14833, n14830, n_13442);
  not g28018 (n_13443, n14832);
  not g28019 (n_13444, n14833);
  and g28020 (n14834, n_13443, n_13444);
  not g28021 (n_13445, n14834);
  and g28022 (n14835, n14781, n_13445);
  not g28023 (n_13446, n14835);
  and g28024 (n14836, n14781, n_13446);
  and g28025 (n14837, n_13445, n_13446);
  not g28026 (n_13447, n14836);
  not g28027 (n_13448, n14837);
  and g28028 (n14838, n_13447, n_13448);
  not g28029 (n_13449, n14685);
  not g28030 (n_13450, n14838);
  and g28031 (n14839, n_13449, n_13450);
  not g28032 (n_13451, n14839);
  and g28033 (n14840, n_13449, n_13451);
  and g28034 (n14841, n_13450, n_13451);
  not g28035 (n_13452, n14840);
  not g28036 (n_13453, n14841);
  and g28037 (n14842, n_13452, n_13453);
  and g28038 (n14843, n_13269, n_13289);
  and g28039 (n14844, n_13238, n_13242);
  and g28040 (n14845, n_13275, n_13279);
  and g28041 (n14846, n14844, n14845);
  not g28042 (n_13454, n14844);
  not g28043 (n_13455, n14845);
  and g28044 (n14847, n_13454, n_13455);
  not g28045 (n_13456, n14846);
  not g28046 (n_13457, n14847);
  and g28047 (n14848, n_13456, n_13457);
  and g28048 (n14849, n_13133, n_13142);
  not g28049 (n_13458, n14848);
  and g28050 (n14850, n_13458, n14849);
  not g28051 (n_13459, n14849);
  and g28052 (n14851, n14848, n_13459);
  not g28053 (n_13460, n14850);
  not g28054 (n_13461, n14851);
  and g28055 (n14852, n_13460, n_13461);
  and g28056 (n14853, n_13148, n_13152);
  not g28057 (n_13462, n14852);
  and g28058 (n14854, n_13462, n14853);
  not g28059 (n_13463, n14853);
  and g28060 (n14855, n14852, n_13463);
  not g28061 (n_13464, n14854);
  not g28062 (n_13465, n14855);
  and g28063 (n14856, n_13464, n_13465);
  and g28064 (n14857, n_13231, n_13232);
  not g28065 (n_13466, n14857);
  and g28066 (n14858, n_13252, n_13466);
  not g28067 (n_13467, n14858);
  and g28068 (n14859, n14856, n_13467);
  not g28069 (n_13468, n14856);
  and g28070 (n14860, n_13468, n14858);
  not g28071 (n_13469, n14859);
  not g28072 (n_13470, n14860);
  and g28073 (n14861, n_13469, n_13470);
  not g28074 (n_13471, n14861);
  and g28075 (n14862, n14843, n_13471);
  not g28076 (n_13472, n14843);
  and g28077 (n14863, n_13472, n14861);
  not g28078 (n_13473, n14862);
  not g28079 (n_13474, n14863);
  and g28080 (n14864, n_13473, n_13474);
  and g28081 (n14865, n_13156, n_13259);
  not g28082 (n_13475, n14865);
  and g28083 (n14866, n14864, n_13475);
  not g28084 (n_13476, n14864);
  and g28085 (n14867, n_13476, n14865);
  not g28086 (n_13477, n14866);
  not g28087 (n_13478, n14867);
  and g28088 (n14868, n_13477, n_13478);
  not g28089 (n_13479, n14842);
  not g28090 (n_13480, n14868);
  and g28091 (n14869, n_13479, n_13480);
  and g28092 (n14870, n14842, n14868);
  not g28093 (n_13481, n14869);
  not g28094 (n_13482, n14870);
  and g28095 (n14871, n_13481, n_13482);
  not g28096 (n_13483, n14684);
  not g28097 (n_13484, n14871);
  and g28098 (n14872, n_13483, n_13484);
  and g28099 (n14873, n14684, n14871);
  not g28100 (n_13485, n14872);
  not g28101 (n_13486, n14873);
  and g28102 (n14874, n_13485, n_13486);
  not g28103 (n_13487, n14683);
  not g28104 (n_13488, n14874);
  and g28105 (n14875, n_13487, n_13488);
  and g28106 (n14876, n14683, n14874);
  or g28107 (\asquared[86] , n14875, n14876);
  and g28108 (n14878, n_13487, n_13486);
  not g28109 (n_13489, n14878);
  and g28110 (n14879, n_13485, n_13489);
  and g28111 (n14880, n_13479, n14868);
  not g28112 (n_13490, n14880);
  and g28113 (n14881, n_13451, n_13490);
  and g28114 (n14882, n_13474, n_13477);
  and g28115 (n14883, n_13402, n_13414);
  and g28116 (n14884, n_13328, n_13343);
  and g28117 (n14885, n14883, n14884);
  not g28118 (n_13491, n14883);
  not g28119 (n_13492, n14884);
  and g28120 (n14886, n_13491, n_13492);
  not g28121 (n_13493, n14885);
  not g28122 (n_13494, n14886);
  and g28123 (n14887, n_13493, n_13494);
  and g28124 (n14888, n_13365, n_13380);
  not g28125 (n_13495, n14887);
  and g28126 (n14889, n_13495, n14888);
  not g28127 (n_13496, n14888);
  and g28128 (n14890, n14887, n_13496);
  not g28129 (n_13497, n14889);
  not g28130 (n_13498, n14890);
  and g28131 (n14891, n_13497, n_13498);
  and g28132 (n14892, n_13457, n_13461);
  and g28133 (n14893, n14722, n14765);
  not g28134 (n_13499, n14722);
  not g28135 (n_13500, n14765);
  and g28136 (n14894, n_13499, n_13500);
  not g28137 (n_13501, n14893);
  not g28138 (n_13502, n14894);
  and g28139 (n14895, n_13501, n_13502);
  not g28140 (n_13503, n14895);
  and g28141 (n14896, n14751, n_13503);
  not g28142 (n_13504, n14751);
  and g28143 (n14897, n_13504, n14895);
  not g28144 (n_13505, n14896);
  not g28145 (n_13506, n14897);
  and g28146 (n14898, n_13505, n_13506);
  and g28147 (n14899, n14705, n14800);
  not g28148 (n_13507, n14705);
  not g28149 (n_13508, n14800);
  and g28150 (n14900, n_13507, n_13508);
  not g28151 (n_13509, n14899);
  not g28152 (n_13510, n14900);
  and g28153 (n14901, n_13509, n_13510);
  not g28154 (n_13511, n14901);
  and g28155 (n14902, n14693, n_13511);
  not g28156 (n_13512, n14693);
  and g28157 (n14903, n_13512, n14901);
  not g28158 (n_13513, n14902);
  not g28159 (n_13514, n14903);
  and g28160 (n14904, n_13513, n_13514);
  and g28161 (n14905, n14898, n14904);
  not g28162 (n_13515, n14898);
  not g28163 (n_13516, n14904);
  and g28164 (n14906, n_13515, n_13516);
  not g28165 (n_13517, n14905);
  not g28166 (n_13518, n14906);
  and g28167 (n14907, n_13517, n_13518);
  not g28168 (n_13519, n14892);
  and g28169 (n14908, n_13519, n14907);
  not g28170 (n_13520, n14907);
  and g28171 (n14909, n14892, n_13520);
  not g28172 (n_13521, n14908);
  not g28173 (n_13522, n14909);
  and g28174 (n14910, n_13521, n_13522);
  and g28175 (n14911, n14891, n14910);
  not g28176 (n_13523, n14891);
  not g28177 (n_13524, n14910);
  and g28178 (n14912, n_13523, n_13524);
  not g28179 (n_13525, n14911);
  not g28180 (n_13526, n14912);
  and g28181 (n14913, n_13525, n_13526);
  and g28182 (n14914, n_13436, n_13439);
  and g28183 (n14915, \a[36] , \a[50] );
  and g28184 (n14916, \a[37] , \a[49] );
  not g28185 (n_13527, n14915);
  not g28186 (n_13528, n14916);
  and g28187 (n14917, n_13527, n_13528);
  and g28188 (n14918, n3687, n6325);
  not g28189 (n_13529, n14918);
  not g28191 (n_13530, n14917);
  not g28194 (n_13531, n14921);
  and g28195 (n14922, n_13529, n_13531);
  and g28196 (n14923, n_13530, n14922);
  and g28197 (n14924, \a[63] , n_13531);
  and g28198 (n14925, \a[23] , n14924);
  not g28199 (n_13532, n14923);
  not g28200 (n_13533, n14925);
  and g28201 (n14926, n_13532, n_13533);
  and g28202 (n14927, n3319, n6968);
  and g28203 (n14928, n2972, n7232);
  and g28204 (n14929, n4150, n7433);
  not g28205 (n_13534, n14928);
  not g28206 (n_13535, n14929);
  and g28207 (n14930, n_13534, n_13535);
  not g28208 (n_13536, n14927);
  not g28209 (n_13537, n14930);
  and g28210 (n14931, n_13536, n_13537);
  not g28211 (n_13538, n14931);
  and g28212 (n14932, \a[53] , n_13538);
  and g28213 (n14933, \a[33] , n14932);
  and g28214 (n14934, n_13536, n_13538);
  and g28215 (n14935, \a[34] , \a[52] );
  and g28216 (n14936, \a[35] , \a[51] );
  not g28217 (n_13539, n14935);
  not g28218 (n_13540, n14936);
  and g28219 (n14937, n_13539, n_13540);
  not g28220 (n_13541, n14937);
  and g28221 (n14938, n14934, n_13541);
  not g28222 (n_13542, n14933);
  not g28223 (n_13543, n14938);
  and g28224 (n14939, n_13542, n_13543);
  not g28225 (n_13544, n14926);
  not g28226 (n_13545, n14939);
  and g28227 (n14940, n_13544, n_13545);
  not g28228 (n_13546, n14940);
  and g28229 (n14941, n_13544, n_13546);
  and g28230 (n14942, n_13545, n_13546);
  not g28231 (n_13547, n14941);
  not g28232 (n_13548, n14942);
  and g28233 (n14943, n_13547, n_13548);
  not g28234 (n_13549, n12323);
  not g28235 (n_13550, n14331);
  and g28236 (n14944, n_13549, n_13550);
  and g28237 (n14945, n3452, n11718);
  not g28238 (n_13551, n14945);
  and g28239 (n14946, n6942, n_13551);
  not g28240 (n_13552, n14944);
  and g28241 (n14947, n_13552, n14946);
  not g28242 (n_13553, n14947);
  and g28243 (n14948, n6942, n_13553);
  and g28244 (n14949, n_13551, n_13553);
  and g28245 (n14950, n_13552, n14949);
  not g28246 (n_13554, n14948);
  not g28247 (n_13555, n14950);
  and g28248 (n14951, n_13554, n_13555);
  not g28249 (n_13556, n14943);
  not g28250 (n_13557, n14951);
  and g28251 (n14952, n_13556, n_13557);
  not g28252 (n_13558, n14952);
  and g28253 (n14953, n_13556, n_13558);
  and g28254 (n14954, n_13557, n_13558);
  not g28255 (n_13559, n14953);
  not g28256 (n_13560, n14954);
  and g28257 (n14955, n_13559, n_13560);
  and g28258 (n14956, n2331, n8987);
  and g28259 (n14957, n2800, n10089);
  and g28260 (n14958, n2227, n9509);
  not g28261 (n_13561, n14957);
  not g28262 (n_13562, n14958);
  and g28263 (n14959, n_13561, n_13562);
  not g28264 (n_13563, n14956);
  not g28265 (n_13564, n14959);
  and g28266 (n14960, n_13563, n_13564);
  not g28267 (n_13565, n14960);
  and g28268 (n14961, n_13563, n_13565);
  and g28269 (n14962, \a[27] , \a[59] );
  and g28270 (n14963, \a[28] , \a[58] );
  not g28271 (n_13566, n14962);
  not g28272 (n_13567, n14963);
  and g28273 (n14964, n_13566, n_13567);
  not g28274 (n_13568, n14964);
  and g28275 (n14965, n14961, n_13568);
  and g28276 (n14966, \a[60] , n_13565);
  and g28277 (n14967, \a[26] , n14966);
  not g28278 (n_13569, n14965);
  not g28279 (n_13570, n14967);
  and g28280 (n14968, n_13569, n_13570);
  and g28281 (n14969, \a[32] , \a[54] );
  and g28282 (n14970, n4639, n14969);
  and g28283 (n14971, n4809, n14969);
  and g28284 (n14972, n5344, n5713);
  not g28285 (n_13571, n14971);
  not g28286 (n_13572, n14972);
  and g28287 (n14973, n_13571, n_13572);
  not g28288 (n_13573, n14970);
  not g28289 (n_13574, n14973);
  and g28290 (n14974, n_13573, n_13574);
  not g28291 (n_13575, n14974);
  and g28292 (n14975, n4809, n_13575);
  and g28293 (n14976, n_13573, n_13575);
  not g28294 (n_13576, n4639);
  not g28295 (n_13577, n14969);
  and g28296 (n14977, n_13576, n_13577);
  not g28297 (n_13578, n14977);
  and g28298 (n14978, n14976, n_13578);
  not g28299 (n_13579, n14975);
  not g28300 (n_13580, n14978);
  and g28301 (n14979, n_13579, n_13580);
  not g28302 (n_13581, n14968);
  not g28303 (n_13582, n14979);
  and g28304 (n14980, n_13581, n_13582);
  not g28305 (n_13583, n14980);
  and g28306 (n14981, n_13581, n_13583);
  and g28307 (n14982, n_13582, n_13583);
  not g28308 (n_13584, n14981);
  not g28309 (n_13585, n14982);
  and g28310 (n14983, n_13584, n_13585);
  and g28311 (n14984, \a[39] , \a[47] );
  not g28312 (n_13586, n7073);
  not g28313 (n_13587, n14984);
  and g28314 (n14985, n_13586, n_13587);
  and g28315 (n14986, n4171, n5666);
  not g28316 (n_13588, n14986);
  not g28319 (n_13589, n14985);
  not g28321 (n_13590, n14989);
  and g28322 (n14990, \a[56] , n_13590);
  and g28323 (n14991, \a[30] , n14990);
  and g28324 (n14992, n_13588, n_13590);
  and g28325 (n14993, n_13589, n14992);
  not g28326 (n_13591, n14991);
  not g28327 (n_13592, n14993);
  and g28328 (n14994, n_13591, n_13592);
  not g28329 (n_13593, n14983);
  not g28330 (n_13594, n14994);
  and g28331 (n14995, n_13593, n_13594);
  not g28332 (n_13595, n14995);
  and g28333 (n14996, n_13593, n_13595);
  and g28334 (n14997, n_13594, n_13595);
  not g28335 (n_13596, n14996);
  not g28336 (n_13597, n14997);
  and g28337 (n14998, n_13596, n_13597);
  and g28338 (n14999, n14955, n14998);
  not g28339 (n_13598, n14955);
  not g28340 (n_13599, n14998);
  and g28341 (n15000, n_13598, n_13599);
  not g28342 (n_13600, n14999);
  not g28343 (n_13601, n15000);
  and g28344 (n15001, n_13600, n_13601);
  not g28345 (n_13602, n14914);
  and g28346 (n15002, n_13602, n15001);
  not g28347 (n_13603, n15001);
  and g28348 (n15003, n14914, n_13603);
  not g28349 (n_13604, n15002);
  not g28350 (n_13605, n15003);
  and g28351 (n15004, n_13604, n_13605);
  and g28352 (n15005, n14913, n15004);
  not g28353 (n_13606, n14913);
  not g28354 (n_13607, n15004);
  and g28355 (n15006, n_13606, n_13607);
  not g28356 (n_13608, n15005);
  not g28357 (n_13609, n15006);
  and g28358 (n15007, n_13608, n_13609);
  not g28359 (n_13610, n14882);
  and g28360 (n15008, n_13610, n15007);
  not g28361 (n_13611, n15008);
  and g28362 (n15009, n_13610, n_13611);
  and g28363 (n15010, n15007, n_13611);
  not g28364 (n_13612, n15009);
  not g28365 (n_13613, n15010);
  and g28366 (n15011, n_13612, n_13613);
  and g28367 (n15012, n_13442, n_13446);
  and g28368 (n15013, n_13465, n_13469);
  and g28369 (n15014, n15012, n15013);
  not g28370 (n_13614, n15012);
  not g28371 (n_13615, n15013);
  and g28372 (n15015, n_13614, n_13615);
  not g28373 (n_13616, n15014);
  not g28374 (n_13617, n15015);
  and g28375 (n15016, n_13616, n_13617);
  and g28376 (n15017, n1904, n9721);
  not g28377 (n_13618, n15017);
  and g28378 (n15018, \a[61] , n_13618);
  and g28379 (n15019, \a[25] , n15018);
  and g28380 (n15020, \a[62] , n_13618);
  and g28381 (n15021, \a[24] , n15020);
  not g28382 (n_13619, n15019);
  not g28383 (n_13620, n15021);
  and g28384 (n15022, n_13619, n_13620);
  not g28385 (n_13621, n14735);
  not g28386 (n_13622, n15022);
  and g28387 (n15023, n_13621, n_13622);
  not g28388 (n_13623, n15023);
  and g28389 (n15024, n_13621, n_13623);
  and g28390 (n15025, n_13622, n_13623);
  not g28391 (n_13624, n15024);
  not g28392 (n_13625, n15025);
  and g28393 (n15026, n_13624, n_13625);
  and g28394 (n15027, n_13393, n_13398);
  and g28395 (n15028, n15026, n15027);
  not g28396 (n_13626, n15026);
  not g28397 (n_13627, n15027);
  and g28398 (n15029, n_13626, n_13627);
  not g28399 (n_13628, n15028);
  not g28400 (n_13629, n15029);
  and g28401 (n15030, n_13628, n_13629);
  and g28402 (n15031, n_13428, n_13432);
  not g28403 (n_13630, n15030);
  and g28404 (n15032, n_13630, n15031);
  not g28405 (n_13631, n15031);
  and g28406 (n15033, n15030, n_13631);
  not g28407 (n_13632, n15032);
  not g28408 (n_13633, n15033);
  and g28409 (n15034, n_13632, n_13633);
  not g28410 (n_13634, n14814);
  and g28411 (n15035, n_13634, n15034);
  not g28412 (n_13635, n15034);
  and g28413 (n15036, n14814, n_13635);
  not g28414 (n_13636, n15035);
  not g28415 (n_13637, n15036);
  and g28416 (n15037, n_13636, n_13637);
  and g28417 (n15038, n_13383, n_13384);
  not g28418 (n_13638, n15038);
  and g28419 (n15039, n_13390, n_13638);
  not g28420 (n_13639, n15039);
  and g28421 (n15040, n15037, n_13639);
  not g28422 (n_13640, n15037);
  and g28423 (n15041, n_13640, n15039);
  not g28424 (n_13641, n15040);
  not g28425 (n_13642, n15041);
  and g28426 (n15042, n_13641, n_13642);
  and g28427 (n15043, n15016, n15042);
  not g28428 (n_13643, n15016);
  not g28429 (n_13644, n15042);
  and g28430 (n15044, n_13643, n_13644);
  not g28431 (n_13645, n15043);
  not g28432 (n_13646, n15044);
  and g28433 (n15045, n_13645, n_13646);
  not g28434 (n_13647, n15011);
  and g28435 (n15046, n_13647, n15045);
  not g28436 (n_13648, n15045);
  and g28437 (n15047, n_13613, n_13648);
  and g28438 (n15048, n_13612, n15047);
  not g28439 (n_13649, n15046);
  not g28440 (n_13650, n15048);
  and g28441 (n15049, n_13649, n_13650);
  not g28442 (n_13651, n15049);
  and g28443 (n15050, n14881, n_13651);
  not g28444 (n_13652, n14881);
  and g28445 (n15051, n_13652, n15049);
  not g28446 (n_13653, n15050);
  not g28447 (n_13654, n15051);
  and g28448 (n15052, n_13653, n_13654);
  not g28449 (n_13655, n15052);
  and g28450 (n15053, n14879, n_13655);
  not g28451 (n_13656, n14879);
  and g28452 (n15054, n_13656, n_13653);
  and g28453 (n15055, n_13654, n15054);
  not g28454 (n_13657, n15053);
  not g28455 (n_13658, n15055);
  and g28456 (\asquared[87] , n_13657, n_13658);
  not g28457 (n_13659, n15054);
  and g28458 (n15057, n_13654, n_13659);
  and g28459 (n15058, n_13611, n_13649);
  and g28460 (n15059, n_13601, n_13604);
  and g28461 (n15060, n_13502, n_13506);
  and g28462 (n15061, n_13546, n_13558);
  and g28463 (n15062, n15060, n15061);
  not g28464 (n_13660, n15060);
  not g28465 (n_13661, n15061);
  and g28466 (n15063, n_13660, n_13661);
  not g28467 (n_13662, n15062);
  not g28468 (n_13663, n15063);
  and g28469 (n15064, n_13662, n_13663);
  and g28470 (n15065, n_13583, n_13595);
  not g28471 (n_13664, n15064);
  and g28472 (n15066, n_13664, n15065);
  not g28473 (n_13665, n15065);
  and g28474 (n15067, n15064, n_13665);
  not g28475 (n_13666, n15066);
  not g28476 (n_13667, n15067);
  and g28477 (n15068, n_13666, n_13667);
  not g28478 (n_13668, n15059);
  and g28479 (n15069, n_13668, n15068);
  not g28480 (n_13669, n15068);
  and g28481 (n15070, n15059, n_13669);
  not g28482 (n_13670, n15069);
  not g28483 (n_13671, n15070);
  and g28484 (n15071, n_13670, n_13671);
  and g28485 (n15072, n_13636, n_13641);
  not g28486 (n_13672, n15071);
  and g28487 (n15073, n_13672, n15072);
  not g28488 (n_13673, n15072);
  and g28489 (n15074, n15071, n_13673);
  not g28490 (n_13674, n15073);
  not g28491 (n_13675, n15074);
  and g28492 (n15075, n_13674, n_13675);
  and g28493 (n15076, n_13617, n_13645);
  not g28494 (n_13676, n15075);
  and g28495 (n15077, n_13676, n15076);
  not g28496 (n_13677, n15076);
  and g28497 (n15078, n15075, n_13677);
  not g28498 (n_13678, n15077);
  not g28499 (n_13679, n15078);
  and g28500 (n15079, n_13678, n_13679);
  and g28501 (n15080, n_13517, n_13521);
  and g28502 (n15081, n_13494, n_13498);
  and g28503 (n15082, n15080, n15081);
  not g28504 (n_13680, n15080);
  not g28505 (n_13681, n15081);
  and g28506 (n15083, n_13680, n_13681);
  not g28507 (n_13682, n15082);
  not g28508 (n_13683, n15083);
  and g28509 (n15084, n_13682, n_13683);
  and g28510 (n15085, n_13629, n_13633);
  and g28511 (n15086, n14976, n14992);
  not g28512 (n_13684, n14976);
  not g28513 (n_13685, n14992);
  and g28514 (n15087, n_13684, n_13685);
  not g28515 (n_13686, n15086);
  not g28516 (n_13687, n15087);
  and g28517 (n15088, n_13686, n_13687);
  not g28518 (n_13688, n15088);
  and g28519 (n15089, n14949, n_13688);
  not g28520 (n_13689, n14949);
  and g28521 (n15090, n_13689, n15088);
  not g28522 (n_13690, n15089);
  not g28523 (n_13691, n15090);
  and g28524 (n15091, n_13690, n_13691);
  and g28525 (n15092, n14934, n14961);
  not g28526 (n_13692, n14934);
  not g28527 (n_13693, n14961);
  and g28528 (n15093, n_13692, n_13693);
  not g28529 (n_13694, n15092);
  not g28530 (n_13695, n15093);
  and g28531 (n15094, n_13694, n_13695);
  not g28532 (n_13696, n15094);
  and g28533 (n15095, n14922, n_13696);
  not g28534 (n_13697, n14922);
  and g28535 (n15096, n_13697, n15094);
  not g28536 (n_13698, n15095);
  not g28537 (n_13699, n15096);
  and g28538 (n15097, n_13698, n_13699);
  not g28539 (n_13700, n15091);
  not g28540 (n_13701, n15097);
  and g28541 (n15098, n_13700, n_13701);
  and g28542 (n15099, n15091, n15097);
  not g28543 (n_13702, n15098);
  not g28544 (n_13703, n15099);
  and g28545 (n15100, n_13702, n_13703);
  not g28546 (n_13704, n15085);
  and g28547 (n15101, n_13704, n15100);
  not g28548 (n_13705, n15100);
  and g28549 (n15102, n15085, n_13705);
  not g28550 (n_13706, n15101);
  not g28551 (n_13707, n15102);
  and g28552 (n15103, n_13706, n_13707);
  and g28553 (n15104, n15084, n15103);
  not g28554 (n_13708, n15084);
  not g28555 (n_13709, n15103);
  and g28556 (n15105, n_13708, n_13709);
  and g28557 (n15106, n_13525, n_13608);
  and g28558 (n15107, \a[44] , \a[62] );
  and g28559 (n15108, \a[25] , n15107);
  not g28560 (n_13710, n15108);
  and g28561 (n15109, n5296, n_13710);
  not g28562 (n_13711, n15109);
  and g28563 (n15110, n_13710, n_13711);
  and g28564 (n15111, \a[25] , \a[62] );
  not g28565 (n_13712, \a[44] );
  not g28566 (n_13713, n15111);
  and g28567 (n15112, n_13712, n_13713);
  not g28568 (n_13714, n15112);
  and g28569 (n15113, n15110, n_13714);
  and g28570 (n15114, n5296, n_13711);
  not g28571 (n_13715, n15113);
  not g28572 (n_13716, n15114);
  and g28573 (n15115, n_13715, n_13716);
  and g28574 (n15116, \a[31] , \a[56] );
  and g28575 (n15117, \a[33] , \a[54] );
  not g28576 (n_13717, n15116);
  not g28577 (n_13718, n15117);
  and g28578 (n15118, n_13717, n_13718);
  and g28579 (n15119, n2598, n7421);
  not g28580 (n_13719, n15119);
  not g28583 (n_13720, n15118);
  not g28585 (n_13721, n15122);
  and g28586 (n15123, \a[47] , n_13721);
  and g28587 (n15124, \a[40] , n15123);
  and g28588 (n15125, n_13719, n_13721);
  and g28589 (n15126, n_13720, n15125);
  not g28590 (n_13722, n15124);
  not g28591 (n_13723, n15126);
  and g28592 (n15127, n_13722, n_13723);
  not g28593 (n_13724, n15115);
  not g28594 (n_13725, n15127);
  and g28595 (n15128, n_13724, n_13725);
  not g28596 (n_13726, n15128);
  and g28597 (n15129, n_13724, n_13726);
  and g28598 (n15130, n_13725, n_13726);
  not g28599 (n_13727, n15129);
  not g28600 (n_13728, n15130);
  and g28601 (n15131, n_13727, n_13728);
  and g28602 (n15132, n_13510, n_13514);
  and g28603 (n15133, n15131, n15132);
  not g28604 (n_13729, n15131);
  not g28605 (n_13730, n15132);
  and g28606 (n15134, n_13729, n_13730);
  not g28607 (n_13731, n15133);
  not g28608 (n_13732, n15134);
  and g28609 (n15135, n_13731, n_13732);
  and g28610 (n15136, n2227, n9512);
  and g28611 (n15137, n2301, n9909);
  and g28612 (n15138, n6196, n11634);
  not g28613 (n_13733, n15137);
  not g28614 (n_13734, n15138);
  and g28615 (n15139, n_13733, n_13734);
  not g28616 (n_13735, n15136);
  not g28617 (n_13736, n15139);
  and g28618 (n15140, n_13735, n_13736);
  not g28619 (n_13737, n15140);
  and g28620 (n15141, n_13735, n_13737);
  and g28621 (n15142, \a[26] , \a[61] );
  and g28622 (n15143, \a[27] , \a[60] );
  not g28623 (n_13738, n15142);
  not g28624 (n_13739, n15143);
  and g28625 (n15144, n_13738, n_13739);
  not g28626 (n_13740, n15144);
  and g28627 (n15145, n15141, n_13740);
  and g28628 (n15146, \a[63] , n_13737);
  and g28629 (n15147, \a[24] , n15146);
  not g28630 (n_13741, n15145);
  not g28631 (n_13742, n15147);
  and g28632 (n15148, n_13741, n_13742);
  and g28633 (n15149, n5083, n6256);
  and g28634 (n15150, n5430, n5888);
  and g28635 (n15151, n4565, n6325);
  not g28636 (n_13743, n15150);
  not g28637 (n_13744, n15151);
  and g28638 (n15152, n_13743, n_13744);
  not g28639 (n_13745, n15149);
  not g28640 (n_13746, n15152);
  and g28641 (n15153, n_13745, n_13746);
  not g28642 (n_13747, n15153);
  and g28643 (n15154, \a[50] , n_13747);
  and g28644 (n15155, \a[37] , n15154);
  and g28645 (n15156, \a[38] , \a[49] );
  and g28646 (n15157, \a[39] , \a[48] );
  not g28647 (n_13748, n15156);
  not g28648 (n_13749, n15157);
  and g28649 (n15158, n_13748, n_13749);
  and g28650 (n15159, n_13745, n_13747);
  not g28651 (n_13750, n15158);
  and g28652 (n15160, n_13750, n15159);
  not g28653 (n_13751, n15155);
  not g28654 (n_13752, n15160);
  and g28655 (n15161, n_13751, n_13752);
  not g28656 (n_13753, n15148);
  not g28657 (n_13754, n15161);
  and g28658 (n15162, n_13753, n_13754);
  not g28659 (n_13755, n15162);
  and g28660 (n15163, n_13753, n_13755);
  and g28661 (n15164, n_13754, n_13755);
  not g28662 (n_13756, n15163);
  not g28663 (n_13757, n15164);
  and g28664 (n15165, n_13756, n_13757);
  and g28665 (n15166, \a[41] , \a[46] );
  and g28666 (n15167, \a[42] , \a[45] );
  not g28667 (n_13758, n15166);
  not g28668 (n_13759, n15167);
  and g28669 (n15168, n_13758, n_13759);
  and g28670 (n15169, n5344, n5560);
  not g28671 (n_13760, n15169);
  not g28674 (n_13761, n15168);
  not g28676 (n_13762, n15172);
  and g28677 (n15173, \a[55] , n_13762);
  and g28678 (n15174, \a[32] , n15173);
  and g28679 (n15175, n_13760, n_13762);
  and g28680 (n15176, n_13761, n15175);
  not g28681 (n_13763, n15174);
  not g28682 (n_13764, n15176);
  and g28683 (n15177, n_13763, n_13764);
  not g28684 (n_13765, n15165);
  not g28685 (n_13766, n15177);
  and g28686 (n15178, n_13765, n_13766);
  not g28687 (n_13767, n15178);
  and g28688 (n15179, n_13765, n_13767);
  and g28689 (n15180, n_13766, n_13767);
  not g28690 (n_13768, n15179);
  not g28691 (n_13769, n15180);
  and g28692 (n15181, n_13768, n_13769);
  not g28693 (n_13770, n15135);
  and g28694 (n15182, n_13770, n15181);
  not g28695 (n_13771, n15181);
  and g28696 (n15183, n15135, n_13771);
  not g28697 (n_13772, n15182);
  not g28698 (n_13773, n15183);
  and g28699 (n15184, n_13772, n_13773);
  and g28700 (n15185, \a[34] , \a[53] );
  and g28701 (n15186, n14598, n15185);
  and g28702 (n15187, n3110, n8985);
  and g28703 (n15188, \a[34] , \a[59] );
  and g28704 (n15189, n13942, n15188);
  not g28705 (n_13774, n15187);
  not g28706 (n_13775, n15189);
  and g28707 (n15190, n_13774, n_13775);
  not g28708 (n_13776, n15186);
  not g28709 (n_13777, n15190);
  and g28710 (n15191, n_13776, n_13777);
  not g28711 (n_13778, n15191);
  and g28712 (n15192, \a[59] , n_13778);
  and g28713 (n15193, \a[28] , n15192);
  and g28714 (n15194, n_13776, n_13778);
  not g28715 (n_13779, n14598);
  not g28716 (n_13780, n15185);
  and g28717 (n15195, n_13779, n_13780);
  not g28718 (n_13781, n15195);
  and g28719 (n15196, n15194, n_13781);
  not g28720 (n_13782, n15193);
  not g28721 (n_13783, n15196);
  and g28722 (n15197, n_13782, n_13783);
  and g28723 (n15198, n_13618, n_13623);
  not g28724 (n_13784, n15197);
  and g28725 (n15199, n_13784, n15198);
  not g28726 (n_13785, n15198);
  and g28727 (n15200, n15197, n_13785);
  not g28728 (n_13786, n15199);
  not g28729 (n_13787, n15200);
  and g28730 (n15201, n_13786, n_13787);
  and g28731 (n15202, n3828, n6968);
  and g28732 (n15203, \a[35] , \a[58] );
  and g28733 (n15204, n13943, n15203);
  not g28734 (n_13788, n15202);
  not g28735 (n_13789, n15204);
  and g28736 (n15205, n_13788, n_13789);
  and g28737 (n15206, \a[29] , \a[58] );
  and g28738 (n15207, \a[36] , \a[51] );
  and g28739 (n15208, n15206, n15207);
  not g28740 (n_13790, n15205);
  not g28741 (n_13791, n15208);
  and g28742 (n15209, n_13790, n_13791);
  not g28743 (n_13792, n15209);
  and g28744 (n15210, \a[52] , n_13792);
  and g28745 (n15211, \a[35] , n15210);
  and g28746 (n15212, n_13791, n_13792);
  not g28747 (n_13793, n15206);
  not g28748 (n_13794, n15207);
  and g28749 (n15213, n_13793, n_13794);
  not g28750 (n_13795, n15213);
  and g28751 (n15214, n15212, n_13795);
  not g28752 (n_13796, n15211);
  not g28753 (n_13797, n15214);
  and g28754 (n15215, n_13796, n_13797);
  not g28755 (n_13798, n15201);
  not g28756 (n_13799, n15215);
  and g28757 (n15216, n_13798, n_13799);
  and g28758 (n15217, n15201, n15215);
  not g28759 (n_13800, n15216);
  not g28760 (n_13801, n15217);
  and g28761 (n15218, n_13800, n_13801);
  and g28762 (n15219, n15184, n15218);
  not g28763 (n_13802, n15184);
  not g28764 (n_13803, n15218);
  and g28765 (n15220, n_13802, n_13803);
  not g28766 (n_13804, n15219);
  not g28767 (n_13805, n15220);
  and g28768 (n15221, n_13804, n_13805);
  not g28769 (n_13806, n15106);
  and g28770 (n15222, n_13806, n15221);
  not g28771 (n_13807, n15221);
  and g28772 (n15223, n15106, n_13807);
  not g28773 (n_13808, n15222);
  not g28774 (n_13809, n15223);
  and g28775 (n15224, n_13808, n_13809);
  not g28776 (n_13810, n15105);
  and g28777 (n15225, n_13810, n15224);
  not g28778 (n_13811, n15104);
  and g28779 (n15226, n_13811, n15225);
  not g28780 (n_13812, n15226);
  and g28781 (n15227, n15224, n_13812);
  and g28782 (n15228, n_13810, n_13812);
  and g28783 (n15229, n_13811, n15228);
  not g28784 (n_13813, n15227);
  not g28785 (n_13814, n15229);
  and g28786 (n15230, n_13813, n_13814);
  not g28787 (n_13815, n15079);
  and g28788 (n15231, n_13815, n15230);
  not g28789 (n_13816, n15230);
  and g28790 (n15232, n15079, n_13816);
  not g28791 (n_13817, n15231);
  not g28792 (n_13818, n15232);
  and g28793 (n15233, n_13817, n_13818);
  not g28794 (n_13819, n15233);
  and g28795 (n15234, n15058, n_13819);
  not g28796 (n_13820, n15058);
  and g28797 (n15235, n_13820, n15233);
  not g28798 (n_13821, n15234);
  not g28799 (n_13822, n15235);
  and g28800 (n15236, n_13821, n_13822);
  not g28801 (n_13823, n15057);
  not g28802 (n_13824, n15236);
  and g28803 (n15237, n_13823, n_13824);
  and g28804 (n15238, n15057, n15236);
  or g28805 (\asquared[88] , n15237, n15238);
  and g28806 (n15240, n_13679, n_13818);
  and g28807 (n15241, n_13670, n_13675);
  and g28808 (n15242, n2331, n9512);
  and g28809 (n15243, n2800, n9085);
  and g28810 (n15244, n2227, n9721);
  not g28811 (n_13825, n15243);
  not g28812 (n_13826, n15244);
  and g28813 (n15245, n_13825, n_13826);
  not g28814 (n_13827, n15242);
  not g28815 (n_13828, n15245);
  and g28816 (n15246, n_13827, n_13828);
  not g28817 (n_13829, n15246);
  and g28818 (n15247, n_13827, n_13829);
  and g28819 (n15248, \a[27] , \a[61] );
  and g28820 (n15249, \a[28] , \a[60] );
  not g28821 (n_13830, n15248);
  not g28822 (n_13831, n15249);
  and g28823 (n15250, n_13830, n_13831);
  not g28824 (n_13832, n15250);
  and g28825 (n15251, n15247, n_13832);
  and g28826 (n15252, \a[62] , n_13829);
  and g28827 (n15253, \a[26] , n15252);
  not g28828 (n_13833, n15251);
  not g28829 (n_13834, n15253);
  and g28830 (n15254, n_13833, n_13834);
  and g28831 (n15255, \a[42] , \a[46] );
  and g28832 (n15256, \a[41] , \a[47] );
  not g28833 (n_13835, n15255);
  not g28834 (n_13836, n15256);
  and g28835 (n15257, n_13835, n_13836);
  and g28836 (n15258, n5344, n5666);
  not g28837 (n_13837, n15258);
  not g28840 (n_13838, n15257);
  not g28842 (n_13839, n15261);
  and g28843 (n15262, \a[57] , n_13839);
  and g28844 (n15263, \a[31] , n15262);
  and g28845 (n15264, n_13837, n_13839);
  and g28846 (n15265, n_13838, n15264);
  not g28847 (n_13840, n15263);
  not g28848 (n_13841, n15265);
  and g28849 (n15266, n_13840, n_13841);
  not g28850 (n_13842, n15254);
  not g28851 (n_13843, n15266);
  and g28852 (n15267, n_13842, n_13843);
  not g28853 (n_13844, n15267);
  and g28854 (n15268, n_13842, n_13844);
  and g28855 (n15269, n_13843, n_13844);
  not g28856 (n_13845, n15268);
  not g28857 (n_13846, n15269);
  and g28858 (n15270, n_13845, n_13846);
  and g28859 (n15271, n3687, n6968);
  and g28860 (n15272, n5031, n7232);
  and g28861 (n15273, n3828, n7433);
  not g28862 (n_13847, n15272);
  not g28863 (n_13848, n15273);
  and g28864 (n15274, n_13847, n_13848);
  not g28865 (n_13849, n15271);
  not g28866 (n_13850, n15274);
  and g28867 (n15275, n_13849, n_13850);
  not g28868 (n_13851, n15275);
  and g28869 (n15276, \a[53] , n_13851);
  and g28870 (n15277, \a[35] , n15276);
  and g28871 (n15278, n_13849, n_13851);
  and g28872 (n15279, \a[37] , \a[51] );
  and g28873 (n15280, \a[36] , \a[52] );
  not g28874 (n_13852, n15279);
  not g28875 (n_13853, n15280);
  and g28876 (n15281, n_13852, n_13853);
  not g28877 (n_13854, n15281);
  and g28878 (n15282, n15278, n_13854);
  not g28879 (n_13855, n15277);
  not g28880 (n_13856, n15282);
  and g28881 (n15283, n_13855, n_13856);
  not g28882 (n_13857, n15270);
  not g28883 (n_13858, n15283);
  and g28884 (n15284, n_13857, n_13858);
  not g28885 (n_13859, n15284);
  and g28886 (n15285, n_13857, n_13859);
  and g28887 (n15286, n_13858, n_13859);
  not g28888 (n_13860, n15285);
  not g28889 (n_13861, n15286);
  and g28890 (n15287, n_13860, n_13861);
  and g28891 (n15288, \a[38] , \a[50] );
  and g28892 (n15289, \a[39] , \a[49] );
  not g28893 (n_13862, n15288);
  not g28894 (n_13863, n15289);
  and g28895 (n15290, n_13862, n_13863);
  and g28896 (n15291, n5083, n6325);
  not g28897 (n_13864, n15291);
  not g28900 (n_13865, n15290);
  not g28902 (n_13866, n15294);
  and g28903 (n15295, n_13864, n_13866);
  and g28904 (n15296, n_13865, n15295);
  and g28905 (n15297, \a[59] , n_13866);
  and g28906 (n15298, \a[29] , n15297);
  not g28907 (n_13867, n15296);
  not g28908 (n_13868, n15298);
  and g28909 (n15299, n_13867, n_13868);
  and g28910 (n15300, \a[30] , \a[58] );
  and g28911 (n15301, \a[32] , \a[56] );
  not g28912 (n_13869, n15300);
  not g28913 (n_13870, n15301);
  and g28914 (n15302, n_13869, n_13870);
  and g28915 (n15303, n2488, n7942);
  not g28916 (n_13871, n15303);
  and g28917 (n15304, n7353, n_13871);
  not g28918 (n_13872, n15302);
  and g28919 (n15305, n_13872, n15304);
  not g28920 (n_13873, n15305);
  and g28921 (n15306, n7353, n_13873);
  and g28922 (n15307, n_13871, n_13873);
  and g28923 (n15308, n_13872, n15307);
  not g28924 (n_13874, n15306);
  not g28925 (n_13875, n15308);
  and g28926 (n15309, n_13874, n_13875);
  not g28927 (n_13876, n15299);
  not g28928 (n_13877, n15309);
  and g28929 (n15310, n_13876, n_13877);
  not g28930 (n_13878, n15310);
  and g28931 (n15311, n_13876, n_13878);
  and g28932 (n15312, n_13877, n_13878);
  not g28933 (n_13879, n15311);
  not g28934 (n_13880, n15312);
  and g28935 (n15313, n_13879, n_13880);
  and g28936 (n15314, n_13687, n_13691);
  and g28937 (n15315, n15313, n15314);
  not g28938 (n_13881, n15313);
  not g28939 (n_13882, n15314);
  and g28940 (n15316, n_13881, n_13882);
  not g28941 (n_13883, n15315);
  not g28942 (n_13884, n15316);
  and g28943 (n15317, n_13883, n_13884);
  and g28944 (n15318, \a[25] , \a[63] );
  not g28945 (n_13885, n15110);
  and g28946 (n15319, n_13885, n15318);
  not g28947 (n_13886, n15318);
  and g28948 (n15320, n15110, n_13886);
  not g28949 (n_13887, n15319);
  not g28950 (n_13888, n15320);
  and g28951 (n15321, n_13887, n_13888);
  not g28952 (n_13889, n15321);
  and g28953 (n15322, n15175, n_13889);
  not g28954 (n_13890, n15175);
  and g28955 (n15323, n_13890, n15321);
  not g28956 (n_13891, n15322);
  not g28957 (n_13892, n15323);
  and g28958 (n15324, n_13891, n_13892);
  and g28959 (n15325, n15317, n15324);
  not g28960 (n_13893, n15317);
  not g28961 (n_13894, n15324);
  and g28962 (n15326, n_13893, n_13894);
  not g28963 (n_13895, n15325);
  not g28964 (n_13896, n15326);
  and g28965 (n15327, n_13895, n_13896);
  not g28966 (n_13897, n15287);
  and g28967 (n15328, n_13897, n15327);
  not g28968 (n_13898, n15328);
  and g28969 (n15329, n_13897, n_13898);
  and g28970 (n15330, n15327, n_13898);
  not g28971 (n_13899, n15329);
  not g28972 (n_13900, n15330);
  and g28973 (n15331, n_13899, n_13900);
  not g28974 (n_13901, n15241);
  not g28975 (n_13902, n15331);
  and g28976 (n15332, n_13901, n_13902);
  not g28977 (n_13903, n15332);
  and g28978 (n15333, n_13901, n_13903);
  and g28979 (n15334, n_13902, n_13903);
  not g28980 (n_13904, n15333);
  not g28981 (n_13905, n15334);
  and g28982 (n15335, n_13904, n_13905);
  and g28983 (n15336, n_13703, n_13706);
  and g28984 (n15337, n_13663, n_13667);
  and g28985 (n15338, n15336, n15337);
  not g28986 (n_13906, n15336);
  not g28987 (n_13907, n15337);
  and g28988 (n15339, n_13906, n_13907);
  not g28989 (n_13908, n15338);
  not g28990 (n_13909, n15339);
  and g28991 (n15340, n_13908, n_13909);
  and g28992 (n15341, n15141, n15194);
  not g28993 (n_13910, n15141);
  not g28994 (n_13911, n15194);
  and g28995 (n15342, n_13910, n_13911);
  not g28996 (n_13912, n15341);
  not g28997 (n_13913, n15342);
  and g28998 (n15343, n_13912, n_13913);
  not g28999 (n_13914, n15343);
  and g29000 (n15344, n15159, n_13914);
  not g29001 (n_13915, n15159);
  and g29002 (n15345, n_13915, n15343);
  not g29003 (n_13916, n15344);
  not g29004 (n_13917, n15345);
  and g29005 (n15346, n_13916, n_13917);
  and g29006 (n15347, n15125, n15212);
  not g29007 (n_13918, n15125);
  not g29008 (n_13919, n15212);
  and g29009 (n15348, n_13918, n_13919);
  not g29010 (n_13920, n15347);
  not g29011 (n_13921, n15348);
  and g29012 (n15349, n_13920, n_13921);
  and g29013 (n15350, \a[33] , \a[55] );
  and g29014 (n15351, \a[34] , \a[54] );
  not g29015 (n_13922, n15350);
  not g29016 (n_13923, n15351);
  and g29017 (n15352, n_13922, n_13923);
  and g29018 (n15353, n4150, n7701);
  not g29019 (n_13924, n15353);
  and g29020 (n15354, n4811, n_13924);
  not g29021 (n_13925, n15352);
  and g29022 (n15355, n_13925, n15354);
  not g29023 (n_13926, n15355);
  and g29024 (n15356, n4811, n_13926);
  and g29025 (n15357, n_13924, n_13926);
  and g29026 (n15358, n_13925, n15357);
  not g29027 (n_13927, n15356);
  not g29028 (n_13928, n15358);
  and g29029 (n15359, n_13927, n_13928);
  not g29030 (n_13929, n15359);
  and g29031 (n15360, n15349, n_13929);
  not g29032 (n_13930, n15360);
  and g29033 (n15361, n15349, n_13930);
  and g29034 (n15362, n_13929, n_13930);
  not g29035 (n_13931, n15361);
  not g29036 (n_13932, n15362);
  and g29037 (n15363, n_13931, n_13932);
  and g29038 (n15364, n_13726, n_13732);
  and g29039 (n15365, n15363, n15364);
  not g29040 (n_13933, n15363);
  not g29041 (n_13934, n15364);
  and g29042 (n15366, n_13933, n_13934);
  not g29043 (n_13935, n15365);
  not g29044 (n_13936, n15366);
  and g29045 (n15367, n_13935, n_13936);
  and g29046 (n15368, n15346, n15367);
  not g29047 (n_13937, n15346);
  not g29048 (n_13938, n15367);
  and g29049 (n15369, n_13937, n_13938);
  not g29050 (n_13939, n15368);
  not g29051 (n_13940, n15369);
  and g29052 (n15370, n_13939, n_13940);
  and g29053 (n15371, n15340, n15370);
  not g29054 (n_13941, n15340);
  not g29055 (n_13942, n15370);
  and g29056 (n15372, n_13941, n_13942);
  not g29057 (n_13943, n15371);
  not g29058 (n_13944, n15372);
  and g29059 (n15373, n_13943, n_13944);
  not g29060 (n_13945, n15335);
  not g29061 (n_13946, n15373);
  and g29062 (n15374, n_13945, n_13946);
  and g29063 (n15375, n15335, n15373);
  not g29064 (n_13947, n15374);
  not g29065 (n_13948, n15375);
  and g29066 (n15376, n_13947, n_13948);
  and g29067 (n15377, n_13808, n_13812);
  and g29068 (n15378, n_13683, n_13811);
  and g29069 (n15379, n_13695, n_13699);
  and g29070 (n15380, n_13784, n_13785);
  not g29071 (n_13949, n15380);
  and g29072 (n15381, n_13800, n_13949);
  and g29073 (n15382, n15379, n15381);
  not g29074 (n_13950, n15379);
  not g29075 (n_13951, n15381);
  and g29076 (n15383, n_13950, n_13951);
  not g29077 (n_13952, n15382);
  not g29078 (n_13953, n15383);
  and g29079 (n15384, n_13952, n_13953);
  and g29080 (n15385, n_13755, n_13767);
  not g29081 (n_13954, n15384);
  and g29082 (n15386, n_13954, n15385);
  not g29083 (n_13955, n15385);
  and g29084 (n15387, n15384, n_13955);
  not g29085 (n_13956, n15386);
  not g29086 (n_13957, n15387);
  and g29087 (n15388, n_13956, n_13957);
  and g29088 (n15389, n_13773, n_13804);
  not g29089 (n_13958, n15389);
  and g29090 (n15390, n15388, n_13958);
  not g29091 (n_13959, n15388);
  and g29092 (n15391, n_13959, n15389);
  not g29093 (n_13960, n15390);
  not g29094 (n_13961, n15391);
  and g29095 (n15392, n_13960, n_13961);
  not g29096 (n_13962, n15378);
  and g29097 (n15393, n_13962, n15392);
  not g29098 (n_13963, n15392);
  and g29099 (n15394, n15378, n_13963);
  not g29100 (n_13964, n15393);
  not g29101 (n_13965, n15394);
  and g29102 (n15395, n_13964, n_13965);
  not g29103 (n_13966, n15377);
  and g29104 (n15396, n_13966, n15395);
  not g29105 (n_13967, n15395);
  and g29106 (n15397, n15377, n_13967);
  not g29107 (n_13968, n15396);
  not g29108 (n_13969, n15397);
  and g29109 (n15398, n_13968, n_13969);
  not g29110 (n_13970, n15376);
  and g29111 (n15399, n_13970, n15398);
  not g29112 (n_13971, n15399);
  and g29113 (n15400, n15398, n_13971);
  and g29114 (n15401, n_13970, n_13971);
  not g29115 (n_13972, n15400);
  not g29116 (n_13973, n15401);
  and g29117 (n15402, n_13972, n_13973);
  and g29118 (n15403, n15240, n15402);
  not g29119 (n_13974, n15240);
  not g29120 (n_13975, n15402);
  and g29121 (n15404, n_13974, n_13975);
  not g29122 (n_13976, n15403);
  not g29123 (n_13977, n15404);
  and g29124 (n15405, n_13976, n_13977);
  and g29125 (n15406, n_13823, n_13821);
  not g29126 (n_13978, n15406);
  and g29127 (n15407, n_13822, n_13978);
  not g29128 (n_13979, n15405);
  and g29129 (n15408, n_13979, n15407);
  not g29130 (n_13980, n15407);
  and g29131 (n15409, n15405, n_13980);
  not g29132 (n_13981, n15408);
  not g29133 (n_13982, n15409);
  and g29134 (\asquared[89] , n_13981, n_13982);
  and g29135 (n15411, n_13968, n_13971);
  and g29136 (n15412, n_13960, n_13964);
  and g29137 (n15413, \a[33] , \a[56] );
  and g29138 (n15414, \a[35] , \a[54] );
  not g29139 (n_13983, n15413);
  not g29140 (n_13984, n15414);
  and g29141 (n15415, n_13983, n_13984);
  and g29142 (n15416, n2972, n7421);
  not g29143 (n_13985, n15416);
  not g29146 (n_13986, n15415);
  not g29148 (n_13987, n15419);
  and g29149 (n15420, n_13985, n_13987);
  and g29150 (n15421, n_13986, n15420);
  and g29151 (n15422, \a[48] , n_13987);
  and g29152 (n15423, \a[41] , n15422);
  not g29153 (n_13988, n15421);
  not g29154 (n_13989, n15423);
  and g29155 (n15424, n_13988, n_13989);
  and g29156 (n15425, n4565, n6968);
  and g29157 (n15426, n3530, n7232);
  and g29158 (n15427, n3687, n7433);
  not g29159 (n_13990, n15426);
  not g29160 (n_13991, n15427);
  and g29161 (n15428, n_13990, n_13991);
  not g29162 (n_13992, n15425);
  not g29163 (n_13993, n15428);
  and g29164 (n15429, n_13992, n_13993);
  not g29165 (n_13994, n15429);
  and g29166 (n15430, \a[53] , n_13994);
  and g29167 (n15431, \a[36] , n15430);
  and g29168 (n15432, n_13992, n_13994);
  not g29169 (n_13995, n7536);
  not g29170 (n_13996, n10556);
  and g29171 (n15433, n_13995, n_13996);
  not g29172 (n_13997, n15433);
  and g29173 (n15434, n15432, n_13997);
  not g29174 (n_13998, n15431);
  not g29175 (n_13999, n15434);
  and g29176 (n15435, n_13998, n_13999);
  not g29177 (n_14000, n15424);
  not g29178 (n_14001, n15435);
  and g29179 (n15436, n_14000, n_14001);
  not g29180 (n_14002, n15436);
  and g29181 (n15437, n_14000, n_14002);
  and g29182 (n15438, n_14001, n_14002);
  not g29183 (n_14003, n15437);
  not g29184 (n_14004, n15438);
  and g29185 (n15439, n_14003, n_14004);
  and g29186 (n15440, n3812, n8436);
  and g29187 (n15441, n2488, n8985);
  and g29188 (n15442, n2865, n8987);
  not g29189 (n_14005, n15441);
  not g29190 (n_14006, n15442);
  and g29191 (n15443, n_14005, n_14006);
  not g29192 (n_14007, n15440);
  not g29193 (n_14008, n15443);
  and g29194 (n15444, n_14007, n_14008);
  not g29195 (n_14009, n15444);
  and g29196 (n15445, \a[59] , n_14009);
  and g29197 (n15446, \a[30] , n15445);
  and g29198 (n15447, n_14007, n_14009);
  and g29199 (n15448, \a[31] , \a[58] );
  and g29200 (n15449, \a[32] , \a[57] );
  not g29201 (n_14010, n15448);
  not g29202 (n_14011, n15449);
  and g29203 (n15450, n_14010, n_14011);
  not g29204 (n_14012, n15450);
  and g29205 (n15451, n15447, n_14012);
  not g29206 (n_14013, n15446);
  not g29207 (n_14014, n15451);
  and g29208 (n15452, n_14013, n_14014);
  not g29209 (n_14015, n15439);
  not g29210 (n_14016, n15452);
  and g29211 (n15453, n_14015, n_14016);
  not g29212 (n_14017, n15453);
  and g29213 (n15454, n_14015, n_14017);
  and g29214 (n15455, n_14016, n_14017);
  not g29215 (n_14018, n15454);
  not g29216 (n_14019, n15455);
  and g29217 (n15456, n_14018, n_14019);
  and g29218 (n15457, n15247, n15278);
  not g29219 (n_14020, n15247);
  not g29220 (n_14021, n15278);
  and g29221 (n15458, n_14020, n_14021);
  not g29222 (n_14022, n15457);
  not g29223 (n_14023, n15458);
  and g29224 (n15459, n_14022, n_14023);
  not g29225 (n_14024, n15459);
  and g29226 (n15460, n15307, n_14024);
  not g29227 (n_14025, n15307);
  and g29228 (n15461, n_14025, n15459);
  not g29229 (n_14026, n15460);
  not g29230 (n_14027, n15461);
  and g29231 (n15462, n_14026, n_14027);
  and g29232 (n15463, \a[45] , \a[62] );
  and g29233 (n15464, \a[27] , n15463);
  not g29234 (n_14028, n15464);
  and g29235 (n15465, n5713, n_14028);
  not g29236 (n_14029, n15465);
  and g29237 (n15466, n_14028, n_14029);
  and g29238 (n15467, \a[27] , \a[62] );
  not g29239 (n_14030, \a[45] );
  not g29240 (n_14031, n15467);
  and g29241 (n15468, n_14030, n_14031);
  not g29242 (n_14032, n15468);
  and g29243 (n15469, n15466, n_14032);
  and g29244 (n15470, n5713, n_14029);
  not g29245 (n_14033, n15469);
  not g29246 (n_14034, n15470);
  and g29247 (n15471, n_14033, n_14034);
  and g29248 (n15472, \a[34] , \a[55] );
  and g29249 (n15473, \a[42] , \a[47] );
  and g29250 (n15474, \a[43] , \a[46] );
  not g29251 (n_14035, n15473);
  not g29252 (n_14036, n15474);
  and g29253 (n15475, n_14035, n_14036);
  and g29254 (n15476, n5018, n5666);
  not g29255 (n_14037, n15476);
  and g29256 (n15477, n15472, n_14037);
  not g29257 (n_14038, n15475);
  and g29258 (n15478, n_14038, n15477);
  not g29259 (n_14039, n15478);
  and g29260 (n15479, n15472, n_14039);
  and g29261 (n15480, n_14037, n_14039);
  and g29262 (n15481, n_14038, n15480);
  not g29263 (n_14040, n15479);
  not g29264 (n_14041, n15481);
  and g29265 (n15482, n_14040, n_14041);
  not g29266 (n_14042, n15471);
  not g29267 (n_14043, n15482);
  and g29268 (n15483, n_14042, n_14043);
  not g29269 (n_14044, n15483);
  and g29270 (n15484, n_14042, n_14044);
  and g29271 (n15485, n_14043, n_14044);
  not g29272 (n_14045, n15484);
  not g29273 (n_14046, n15485);
  and g29274 (n15486, n_14045, n_14046);
  and g29275 (n15487, n2334, n9512);
  not g29276 (n_14047, n15487);
  and g29277 (n15488, \a[60] , n_14047);
  and g29278 (n15489, \a[29] , n15488);
  and g29279 (n15490, \a[61] , n_14047);
  and g29280 (n15491, \a[28] , n15490);
  not g29281 (n_14048, n15489);
  not g29282 (n_14049, n15491);
  and g29283 (n15492, n_14048, n_14049);
  not g29284 (n_14050, n15357);
  not g29285 (n_14051, n15492);
  and g29286 (n15493, n_14050, n_14051);
  not g29287 (n_14052, n15493);
  and g29288 (n15494, n_14050, n_14052);
  and g29289 (n15495, n_14051, n_14052);
  not g29290 (n_14053, n15494);
  not g29291 (n_14054, n15495);
  and g29292 (n15496, n_14053, n_14054);
  not g29293 (n_14055, n15486);
  and g29294 (n15497, n_14055, n15496);
  not g29295 (n_14056, n15496);
  and g29296 (n15498, n15486, n_14056);
  not g29297 (n_14057, n15497);
  not g29298 (n_14058, n15498);
  and g29299 (n15499, n_14057, n_14058);
  not g29300 (n_14059, n15499);
  and g29301 (n15500, n15462, n_14059);
  not g29302 (n_14060, n15500);
  and g29303 (n15501, n15462, n_14060);
  and g29304 (n15502, n_14059, n_14060);
  not g29305 (n_14061, n15501);
  not g29306 (n_14062, n15502);
  and g29307 (n15503, n_14061, n_14062);
  not g29308 (n_14063, n15456);
  not g29309 (n_14064, n15503);
  and g29310 (n15504, n_14063, n_14064);
  not g29311 (n_14065, n15504);
  and g29312 (n15505, n_14063, n_14065);
  and g29313 (n15506, n_14064, n_14065);
  not g29314 (n_14066, n15505);
  not g29315 (n_14067, n15506);
  and g29316 (n15507, n_14066, n_14067);
  not g29317 (n_14068, n15412);
  not g29318 (n_14069, n15507);
  and g29319 (n15508, n_14068, n_14069);
  not g29320 (n_14070, n15508);
  and g29321 (n15509, n_14068, n_14070);
  and g29322 (n15510, n_14069, n_14070);
  not g29323 (n_14071, n15509);
  not g29324 (n_14072, n15510);
  and g29325 (n15511, n_14071, n_14072);
  and g29326 (n15512, n_13913, n_13917);
  and g29327 (n15513, n_13887, n_13892);
  and g29328 (n15514, n15512, n15513);
  not g29329 (n_14073, n15512);
  not g29330 (n_14074, n15513);
  and g29331 (n15515, n_14073, n_14074);
  not g29332 (n_14075, n15514);
  not g29333 (n_14076, n15515);
  and g29334 (n15516, n_14075, n_14076);
  and g29335 (n15517, n_13921, n_13930);
  not g29336 (n_14077, n15516);
  and g29337 (n15518, n_14077, n15517);
  not g29338 (n_14078, n15517);
  and g29339 (n15519, n15516, n_14078);
  not g29340 (n_14079, n15518);
  not g29341 (n_14080, n15519);
  and g29342 (n15520, n_14079, n_14080);
  and g29343 (n15521, n_13953, n_13957);
  not g29344 (n_14081, n15520);
  and g29345 (n15522, n_14081, n15521);
  not g29346 (n_14082, n15521);
  and g29347 (n15523, n15520, n_14082);
  not g29348 (n_14083, n15522);
  not g29349 (n_14084, n15523);
  and g29350 (n15524, n_14083, n_14084);
  and g29351 (n15525, n_13936, n_13939);
  not g29352 (n_14085, n15525);
  and g29353 (n15526, n15524, n_14085);
  not g29354 (n_14086, n15524);
  and g29355 (n15527, n_14086, n15525);
  not g29356 (n_14087, n15526);
  not g29357 (n_14088, n15527);
  and g29358 (n15528, n_14087, n_14088);
  not g29359 (n_14089, n15511);
  and g29360 (n15529, n_14089, n15528);
  not g29361 (n_14090, n15529);
  and g29362 (n15530, n_14089, n_14090);
  and g29363 (n15531, n15528, n_14090);
  not g29364 (n_14091, n15530);
  not g29365 (n_14092, n15531);
  and g29366 (n15532, n_14091, n_14092);
  and g29367 (n15533, n_13945, n15373);
  not g29368 (n_14093, n15533);
  and g29369 (n15534, n_13903, n_14093);
  and g29370 (n15535, n_13909, n_13943);
  and g29371 (n15536, n_13895, n_13898);
  and g29372 (n15537, n_13878, n_13884);
  and g29373 (n15538, n_13844, n_13859);
  and g29374 (n15539, n15537, n15538);
  not g29375 (n_14094, n15537);
  not g29376 (n_14095, n15538);
  and g29377 (n15540, n_14094, n_14095);
  not g29378 (n_14096, n15539);
  not g29379 (n_14097, n15540);
  and g29380 (n15541, n_14096, n_14097);
  and g29381 (n15542, n15264, n15295);
  not g29382 (n_14098, n15264);
  not g29383 (n_14099, n15295);
  and g29384 (n15543, n_14098, n_14099);
  not g29385 (n_14100, n15542);
  not g29386 (n_14101, n15543);
  and g29387 (n15544, n_14100, n_14101);
  and g29388 (n15545, \a[39] , \a[50] );
  and g29389 (n15546, \a[40] , \a[49] );
  not g29390 (n_14102, n15545);
  not g29391 (n_14103, n15546);
  and g29392 (n15547, n_14102, n_14103);
  and g29393 (n15548, n4171, n6325);
  not g29394 (n_14104, n15548);
  not g29396 (n_14105, n15547);
  not g29399 (n_14106, n15551);
  and g29400 (n15552, \a[63] , n_14106);
  and g29401 (n15553, \a[26] , n15552);
  and g29402 (n15554, n_14104, n_14106);
  and g29403 (n15555, n_14105, n15554);
  not g29404 (n_14107, n15553);
  not g29405 (n_14108, n15555);
  and g29406 (n15556, n_14107, n_14108);
  not g29407 (n_14109, n15556);
  and g29408 (n15557, n15544, n_14109);
  not g29409 (n_14110, n15557);
  and g29410 (n15558, n15544, n_14110);
  and g29411 (n15559, n_14109, n_14110);
  not g29412 (n_14111, n15558);
  not g29413 (n_14112, n15559);
  and g29414 (n15560, n_14111, n_14112);
  not g29415 (n_14113, n15541);
  and g29416 (n15561, n_14113, n15560);
  not g29417 (n_14114, n15560);
  and g29418 (n15562, n15541, n_14114);
  not g29419 (n_14115, n15561);
  not g29420 (n_14116, n15562);
  and g29421 (n15563, n_14115, n_14116);
  not g29422 (n_14117, n15536);
  and g29423 (n15564, n_14117, n15563);
  not g29424 (n_14118, n15563);
  and g29425 (n15565, n15536, n_14118);
  not g29426 (n_14119, n15564);
  not g29427 (n_14120, n15565);
  and g29428 (n15566, n_14119, n_14120);
  not g29429 (n_14121, n15535);
  and g29430 (n15567, n_14121, n15566);
  not g29431 (n_14122, n15566);
  and g29432 (n15568, n15535, n_14122);
  not g29433 (n_14123, n15567);
  not g29434 (n_14124, n15568);
  and g29435 (n15569, n_14123, n_14124);
  not g29436 (n_14125, n15534);
  and g29437 (n15570, n_14125, n15569);
  not g29438 (n_14126, n15570);
  and g29439 (n15571, n15569, n_14126);
  and g29440 (n15572, n_14125, n_14126);
  not g29441 (n_14127, n15571);
  not g29442 (n_14128, n15572);
  and g29443 (n15573, n_14127, n_14128);
  not g29444 (n_14129, n15532);
  not g29445 (n_14130, n15573);
  and g29446 (n15574, n_14129, n_14130);
  and g29447 (n15575, n15532, n_14128);
  and g29448 (n15576, n_14127, n15575);
  not g29449 (n_14131, n15574);
  not g29450 (n_14132, n15576);
  and g29451 (n15577, n_14131, n_14132);
  not g29452 (n_14133, n15411);
  and g29453 (n15578, n_14133, n15577);
  not g29454 (n_14134, n15577);
  and g29455 (n15579, n15411, n_14134);
  not g29456 (n_14135, n15578);
  not g29457 (n_14136, n15579);
  and g29458 (n15580, n_14135, n_14136);
  and g29459 (n15581, n_13976, n_13980);
  not g29460 (n_14137, n15581);
  and g29461 (n15582, n_13977, n_14137);
  not g29462 (n_14138, n15580);
  and g29463 (n15583, n_14138, n15582);
  not g29464 (n_14139, n15582);
  and g29465 (n15584, n15580, n_14139);
  not g29466 (n_14140, n15583);
  not g29467 (n_14141, n15584);
  and g29468 (\asquared[90] , n_14140, n_14141);
  and g29469 (n15586, n_14136, n_14139);
  not g29470 (n_14142, n15586);
  and g29471 (n15587, n_14135, n_14142);
  and g29472 (n15588, n_14126, n_14131);
  and g29473 (n15589, n_14084, n_14087);
  and g29474 (n15590, n_14060, n_14065);
  and g29475 (n15591, n15466, n15480);
  not g29476 (n_14143, n15466);
  not g29477 (n_14144, n15480);
  and g29478 (n15592, n_14143, n_14144);
  not g29479 (n_14145, n15591);
  not g29480 (n_14146, n15592);
  and g29481 (n15593, n_14145, n_14146);
  not g29482 (n_14147, n15593);
  and g29483 (n15594, n15420, n_14147);
  not g29484 (n_14148, n15420);
  and g29485 (n15595, n_14148, n15593);
  not g29486 (n_14149, n15594);
  not g29487 (n_14150, n15595);
  and g29488 (n15596, n_14149, n_14150);
  and g29489 (n15597, n_14055, n_14056);
  not g29490 (n_14151, n15597);
  and g29491 (n15598, n_14044, n_14151);
  and g29492 (n15599, n_14002, n_14017);
  and g29493 (n15600, n15598, n15599);
  not g29494 (n_14152, n15598);
  not g29495 (n_14153, n15599);
  and g29496 (n15601, n_14152, n_14153);
  not g29497 (n_14154, n15600);
  not g29498 (n_14155, n15601);
  and g29499 (n15602, n_14154, n_14155);
  and g29500 (n15603, n15596, n15602);
  not g29501 (n_14156, n15596);
  not g29502 (n_14157, n15602);
  and g29503 (n15604, n_14156, n_14157);
  not g29504 (n_14158, n15603);
  not g29505 (n_14159, n15604);
  and g29506 (n15605, n_14158, n_14159);
  not g29507 (n_14160, n15590);
  and g29508 (n15606, n_14160, n15605);
  not g29509 (n_14161, n15605);
  and g29510 (n15607, n15590, n_14161);
  not g29511 (n_14162, n15606);
  not g29512 (n_14163, n15607);
  and g29513 (n15608, n_14162, n_14163);
  not g29514 (n_14164, n15608);
  and g29515 (n15609, n15589, n_14164);
  not g29516 (n_14165, n15589);
  and g29517 (n15610, n_14165, n15608);
  not g29518 (n_14166, n15609);
  not g29519 (n_14167, n15610);
  and g29520 (n15611, n_14166, n_14167);
  and g29521 (n15612, n_14070, n_14090);
  not g29522 (n_14168, n15611);
  and g29523 (n15613, n_14168, n15612);
  not g29524 (n_14169, n15612);
  and g29525 (n15614, n15611, n_14169);
  not g29526 (n_14170, n15613);
  not g29527 (n_14171, n15614);
  and g29528 (n15615, n_14170, n_14171);
  and g29529 (n15616, n_14119, n_14123);
  and g29530 (n15617, n15432, n15447);
  not g29531 (n_14172, n15432);
  not g29532 (n_14173, n15447);
  and g29533 (n15618, n_14172, n_14173);
  not g29534 (n_14174, n15617);
  not g29535 (n_14175, n15618);
  and g29536 (n15619, n_14174, n_14175);
  not g29537 (n_14176, n15619);
  and g29538 (n15620, n15554, n_14176);
  not g29539 (n_14177, n15554);
  and g29540 (n15621, n_14177, n15619);
  not g29541 (n_14178, n15620);
  not g29542 (n_14179, n15621);
  and g29543 (n15622, n_14178, n_14179);
  and g29544 (n15623, n_14076, n_14080);
  not g29545 (n_14180, n15622);
  and g29546 (n15624, n_14180, n15623);
  not g29547 (n_14181, n15623);
  and g29548 (n15625, n15622, n_14181);
  not g29549 (n_14182, n15624);
  not g29550 (n_14183, n15625);
  and g29551 (n15626, n_14182, n_14183);
  and g29552 (n15627, \a[33] , \a[57] );
  and g29553 (n15628, \a[34] , \a[56] );
  not g29554 (n_14184, n15627);
  not g29555 (n_14185, n15628);
  and g29556 (n15629, n_14184, n_14185);
  and g29557 (n15630, n4150, n8200);
  and g29558 (n15631, n2972, n11718);
  and g29559 (n15632, n3319, n9161);
  not g29560 (n_14186, n15631);
  not g29561 (n_14187, n15632);
  and g29562 (n15633, n_14186, n_14187);
  not g29563 (n_14188, n15630);
  not g29564 (n_14189, n15633);
  and g29565 (n15634, n_14188, n_14189);
  not g29566 (n_14190, n15634);
  and g29567 (n15635, n_14188, n_14190);
  not g29568 (n_14191, n15629);
  and g29569 (n15636, n_14191, n15635);
  and g29570 (n15637, \a[55] , n_14190);
  and g29571 (n15638, \a[35] , n15637);
  not g29572 (n_14192, n15636);
  not g29573 (n_14193, n15638);
  and g29574 (n15639, n_14192, n_14193);
  and g29575 (n15640, n4565, n7433);
  and g29576 (n15641, n3530, n10905);
  and g29577 (n15642, n3687, n7699);
  not g29578 (n_14194, n15641);
  not g29579 (n_14195, n15642);
  and g29580 (n15643, n_14194, n_14195);
  not g29581 (n_14196, n15640);
  not g29582 (n_14197, n15643);
  and g29583 (n15644, n_14196, n_14197);
  not g29584 (n_14198, n15644);
  and g29585 (n15645, \a[54] , n_14198);
  and g29586 (n15646, \a[36] , n15645);
  and g29587 (n15647, n_14196, n_14198);
  and g29588 (n15648, \a[38] , \a[52] );
  not g29589 (n_14199, n7435);
  not g29590 (n_14200, n15648);
  and g29591 (n15649, n_14199, n_14200);
  not g29592 (n_14201, n15649);
  and g29593 (n15650, n15647, n_14201);
  not g29594 (n_14202, n15646);
  not g29595 (n_14203, n15650);
  and g29596 (n15651, n_14202, n_14203);
  not g29597 (n_14204, n15639);
  not g29598 (n_14205, n15651);
  and g29599 (n15652, n_14204, n_14205);
  not g29600 (n_14206, n15652);
  and g29601 (n15653, n_14204, n_14206);
  and g29602 (n15654, n_14205, n_14206);
  not g29603 (n_14207, n15653);
  not g29604 (n_14208, n15654);
  and g29605 (n15655, n_14207, n_14208);
  and g29606 (n15656, n5296, n5666);
  and g29607 (n15657, n4639, n8578);
  and g29608 (n15658, n5018, n6252);
  not g29609 (n_14209, n15657);
  not g29610 (n_14210, n15658);
  and g29611 (n15659, n_14209, n_14210);
  not g29612 (n_14211, n15656);
  not g29613 (n_14212, n15659);
  and g29614 (n15660, n_14211, n_14212);
  not g29615 (n_14213, n15660);
  and g29616 (n15661, \a[48] , n_14213);
  and g29617 (n15662, \a[42] , n15661);
  and g29618 (n15663, n_14211, n_14213);
  not g29619 (n_14214, n7747);
  not g29620 (n_14215, n8053);
  and g29621 (n15664, n_14214, n_14215);
  not g29622 (n_14216, n15664);
  and g29623 (n15665, n15663, n_14216);
  not g29624 (n_14217, n15662);
  not g29625 (n_14218, n15665);
  and g29626 (n15666, n_14217, n_14218);
  not g29627 (n_14219, n15655);
  not g29628 (n_14220, n15666);
  and g29629 (n15667, n_14219, n_14220);
  not g29630 (n_14221, n15667);
  and g29631 (n15668, n_14219, n_14221);
  and g29632 (n15669, n_14220, n_14221);
  not g29633 (n_14222, n15668);
  not g29634 (n_14223, n15669);
  and g29635 (n15670, n_14222, n_14223);
  not g29636 (n_14224, n15670);
  and g29637 (n15671, n15626, n_14224);
  not g29638 (n_14225, n15626);
  and g29639 (n15672, n_14225, n15670);
  not g29640 (n_14226, n15616);
  not g29641 (n_14227, n15672);
  and g29642 (n15673, n_14226, n_14227);
  not g29643 (n_14228, n15671);
  and g29644 (n15674, n_14228, n15673);
  not g29645 (n_14229, n15674);
  and g29646 (n15675, n_14226, n_14229);
  and g29647 (n15676, n_14227, n_14229);
  and g29648 (n15677, n_14228, n15676);
  not g29649 (n_14230, n15675);
  not g29650 (n_14231, n15677);
  and g29651 (n15678, n_14230, n_14231);
  and g29652 (n15679, n_14097, n_14116);
  and g29653 (n15680, n_14023, n_14027);
  and g29654 (n15681, n5413, n6325);
  and g29655 (n15682, n3984, n9934);
  and g29656 (n15683, n4171, n6564);
  not g29657 (n_14232, n15682);
  not g29658 (n_14233, n15683);
  and g29659 (n15684, n_14232, n_14233);
  not g29660 (n_14234, n15681);
  not g29661 (n_14235, n15684);
  and g29662 (n15685, n_14234, n_14235);
  not g29663 (n_14236, n15685);
  and g29664 (n15686, n7774, n_14236);
  and g29665 (n15687, n_14234, n_14236);
  and g29666 (n15688, \a[41] , \a[49] );
  and g29667 (n15689, \a[40] , \a[50] );
  not g29668 (n_14237, n15688);
  not g29669 (n_14238, n15689);
  and g29670 (n15690, n_14237, n_14238);
  not g29671 (n_14239, n15690);
  and g29672 (n15691, n15687, n_14239);
  not g29673 (n_14240, n15686);
  not g29674 (n_14241, n15691);
  and g29675 (n15692, n_14240, n_14241);
  not g29676 (n_14242, n15680);
  not g29677 (n_14243, n15692);
  and g29678 (n15693, n_14242, n_14243);
  not g29679 (n_14244, n15693);
  and g29680 (n15694, n_14242, n_14244);
  and g29681 (n15695, n_14243, n_14244);
  not g29682 (n_14245, n15694);
  not g29683 (n_14246, n15695);
  and g29684 (n15696, n_14245, n_14246);
  and g29685 (n15697, n_14101, n_14110);
  and g29686 (n15698, n15696, n15697);
  not g29687 (n_14247, n15696);
  not g29688 (n_14248, n15697);
  and g29689 (n15699, n_14247, n_14248);
  not g29690 (n_14249, n15698);
  not g29691 (n_14250, n15699);
  and g29692 (n15700, n_14249, n_14250);
  and g29693 (n15701, n2334, n9721);
  and g29694 (n15702, n2331, n9792);
  and g29695 (n15703, n2041, n9909);
  not g29696 (n_14251, n15702);
  not g29697 (n_14252, n15703);
  and g29698 (n15704, n_14251, n_14252);
  not g29699 (n_14253, n15701);
  not g29700 (n_14254, n15704);
  and g29701 (n15705, n_14253, n_14254);
  not g29702 (n_14255, n15705);
  and g29703 (n15706, n_14253, n_14255);
  and g29704 (n15707, \a[28] , \a[62] );
  and g29705 (n15708, \a[29] , \a[61] );
  not g29706 (n_14256, n15707);
  not g29707 (n_14257, n15708);
  and g29708 (n15709, n_14256, n_14257);
  not g29709 (n_14258, n15709);
  and g29710 (n15710, n15706, n_14258);
  and g29711 (n15711, \a[63] , n_14255);
  and g29712 (n15712, \a[27] , n15711);
  not g29713 (n_14259, n15710);
  not g29714 (n_14260, n15712);
  and g29715 (n15713, n_14259, n_14260);
  and g29716 (n15714, n_14047, n_14052);
  and g29717 (n15715, n3812, n8987);
  and g29718 (n15716, n2488, n10089);
  and g29719 (n15717, n2865, n9509);
  not g29720 (n_14261, n15716);
  not g29721 (n_14262, n15717);
  and g29722 (n15718, n_14261, n_14262);
  not g29723 (n_14263, n15715);
  not g29724 (n_14264, n15718);
  and g29725 (n15719, n_14263, n_14264);
  and g29726 (n15720, \a[31] , \a[59] );
  not g29727 (n_14265, n14420);
  not g29728 (n_14266, n15720);
  and g29729 (n15721, n_14265, n_14266);
  not g29730 (n_14267, n15721);
  and g29731 (n15722, n_14263, n_14267);
  and g29732 (n15723, \a[30] , \a[60] );
  not g29733 (n_14268, n15722);
  not g29734 (n_14269, n15723);
  and g29735 (n15724, n_14268, n_14269);
  not g29736 (n_14270, n15719);
  not g29737 (n_14271, n15724);
  and g29738 (n15725, n_14270, n_14271);
  not g29739 (n_14272, n15714);
  and g29740 (n15726, n_14272, n15725);
  not g29741 (n_14273, n15726);
  and g29742 (n15727, n_14272, n_14273);
  and g29743 (n15728, n15725, n_14273);
  not g29744 (n_14274, n15727);
  not g29745 (n_14275, n15728);
  and g29746 (n15729, n_14274, n_14275);
  not g29747 (n_14276, n15713);
  not g29748 (n_14277, n15729);
  and g29749 (n15730, n_14276, n_14277);
  and g29750 (n15731, n15713, n_14275);
  and g29751 (n15732, n_14274, n15731);
  not g29752 (n_14278, n15730);
  not g29753 (n_14279, n15732);
  and g29754 (n15733, n_14278, n_14279);
  and g29755 (n15734, n15700, n15733);
  not g29756 (n_14280, n15734);
  and g29757 (n15735, n15700, n_14280);
  and g29758 (n15736, n15733, n_14280);
  not g29759 (n_14281, n15735);
  not g29760 (n_14282, n15736);
  and g29761 (n15737, n_14281, n_14282);
  not g29762 (n_14283, n15679);
  not g29763 (n_14284, n15737);
  and g29764 (n15738, n_14283, n_14284);
  not g29765 (n_14285, n15738);
  and g29766 (n15739, n_14283, n_14285);
  and g29767 (n15740, n_14284, n_14285);
  not g29768 (n_14286, n15739);
  not g29769 (n_14287, n15740);
  and g29770 (n15741, n_14286, n_14287);
  not g29771 (n_14288, n15678);
  not g29772 (n_14289, n15741);
  and g29773 (n15742, n_14288, n_14289);
  not g29774 (n_14290, n15742);
  and g29775 (n15743, n_14288, n_14290);
  and g29776 (n15744, n_14289, n_14290);
  not g29777 (n_14291, n15743);
  not g29778 (n_14292, n15744);
  and g29779 (n15745, n_14291, n_14292);
  not g29780 (n_14293, n15615);
  and g29781 (n15746, n_14293, n15745);
  not g29782 (n_14294, n15745);
  and g29783 (n15747, n15615, n_14294);
  not g29784 (n_14295, n15746);
  not g29785 (n_14296, n15747);
  and g29786 (n15748, n_14295, n_14296);
  not g29787 (n_14297, n15748);
  and g29788 (n15749, n15588, n_14297);
  not g29789 (n_14298, n15588);
  and g29790 (n15750, n_14298, n15748);
  not g29791 (n_14299, n15749);
  not g29792 (n_14300, n15750);
  and g29793 (n15751, n_14299, n_14300);
  not g29794 (n_14301, n15751);
  and g29795 (n15752, n15587, n_14301);
  not g29796 (n_14302, n15587);
  and g29797 (n15753, n_14302, n_14299);
  and g29798 (n15754, n_14300, n15753);
  not g29799 (n_14303, n15752);
  not g29800 (n_14304, n15754);
  and g29801 (\asquared[91] , n_14303, n_14304);
  not g29802 (n_14305, n15753);
  and g29803 (n15756, n_14300, n_14305);
  and g29804 (n15757, n_14171, n_14296);
  and g29805 (n15758, n_14146, n_14150);
  and g29806 (n15759, \a[34] , \a[57] );
  and g29807 (n15760, \a[36] , \a[55] );
  not g29808 (n_14306, n15759);
  not g29809 (n_14307, n15760);
  and g29810 (n15761, n_14306, n_14307);
  and g29811 (n15762, n4595, n11718);
  not g29812 (n_14308, n15762);
  and g29813 (n15763, n7972, n_14308);
  not g29814 (n_14309, n15761);
  and g29815 (n15764, n_14309, n15763);
  not g29816 (n_14310, n15764);
  and g29817 (n15765, n7972, n_14310);
  and g29818 (n15766, n_14308, n_14310);
  and g29819 (n15767, n_14309, n15766);
  not g29820 (n_14311, n15765);
  not g29821 (n_14312, n15767);
  and g29822 (n15768, n_14311, n_14312);
  not g29823 (n_14313, n15758);
  not g29824 (n_14314, n15768);
  and g29825 (n15769, n_14313, n_14314);
  not g29826 (n_14315, n15769);
  and g29827 (n15770, n_14313, n_14315);
  and g29828 (n15771, n_14314, n_14315);
  not g29829 (n_14316, n15770);
  not g29830 (n_14317, n15771);
  and g29831 (n15772, n_14316, n_14317);
  and g29832 (n15773, n_14175, n_14179);
  and g29833 (n15774, n15772, n15773);
  not g29834 (n_14318, n15772);
  not g29835 (n_14319, n15773);
  and g29836 (n15775, n_14318, n_14319);
  not g29837 (n_14320, n15774);
  not g29838 (n_14321, n15775);
  and g29839 (n15776, n_14320, n_14321);
  and g29840 (n15777, n_14155, n_14158);
  and g29841 (n15778, n3143, n8987);
  and g29842 (n15779, n2598, n10089);
  and g29843 (n15780, n3812, n9509);
  not g29844 (n_14322, n15779);
  not g29845 (n_14323, n15780);
  and g29846 (n15781, n_14322, n_14323);
  not g29847 (n_14324, n15778);
  not g29848 (n_14325, n15781);
  and g29849 (n15782, n_14324, n_14325);
  not g29850 (n_14326, n15782);
  and g29851 (n15783, n_14324, n_14326);
  and g29852 (n15784, \a[33] , \a[58] );
  not g29853 (n_14327, n8308);
  not g29854 (n_14328, n15784);
  and g29855 (n15785, n_14327, n_14328);
  not g29856 (n_14329, n15785);
  and g29857 (n15786, n15783, n_14329);
  and g29858 (n15787, \a[60] , n_14326);
  and g29859 (n15788, \a[31] , n15787);
  not g29860 (n_14330, n15786);
  not g29861 (n_14331, n15788);
  and g29862 (n15789, n_14330, n_14331);
  and g29863 (n15790, n5083, n7433);
  and g29864 (n15791, n5430, n10905);
  and g29865 (n15792, n4565, n7699);
  not g29866 (n_14332, n15791);
  not g29867 (n_14333, n15792);
  and g29868 (n15793, n_14332, n_14333);
  not g29869 (n_14334, n15790);
  not g29870 (n_14335, n15793);
  and g29871 (n15794, n_14334, n_14335);
  not g29872 (n_14336, n15794);
  and g29873 (n15795, \a[37] , n_14336);
  and g29874 (n15796, \a[54] , n15795);
  and g29875 (n15797, n_14334, n_14336);
  and g29876 (n15798, \a[38] , \a[53] );
  and g29877 (n15799, \a[39] , \a[52] );
  not g29878 (n_14337, n15798);
  not g29879 (n_14338, n15799);
  and g29880 (n15800, n_14337, n_14338);
  not g29881 (n_14339, n15800);
  and g29882 (n15801, n15797, n_14339);
  not g29883 (n_14340, n15796);
  not g29884 (n_14341, n15801);
  and g29885 (n15802, n_14340, n_14341);
  not g29886 (n_14342, n15687);
  not g29887 (n_14343, n15802);
  and g29888 (n15803, n_14342, n_14343);
  not g29889 (n_14344, n15803);
  and g29890 (n15804, n_14342, n_14344);
  and g29891 (n15805, n_14343, n_14344);
  not g29892 (n_14345, n15804);
  not g29893 (n_14346, n15805);
  and g29894 (n15806, n_14345, n_14346);
  not g29895 (n_14347, n15789);
  not g29896 (n_14348, n15806);
  and g29897 (n15807, n_14347, n_14348);
  not g29898 (n_14349, n15807);
  and g29899 (n15808, n_14347, n_14349);
  and g29900 (n15809, n_14348, n_14349);
  not g29901 (n_14350, n15808);
  not g29902 (n_14351, n15809);
  and g29903 (n15810, n_14350, n_14351);
  not g29904 (n_14352, n15777);
  not g29905 (n_14353, n15810);
  and g29906 (n15811, n_14352, n_14353);
  not g29907 (n_14354, n15811);
  and g29908 (n15812, n_14352, n_14354);
  and g29909 (n15813, n_14353, n_14354);
  not g29910 (n_14355, n15812);
  not g29911 (n_14356, n15813);
  and g29912 (n15814, n_14355, n_14356);
  not g29913 (n_14357, n15814);
  and g29914 (n15815, n15776, n_14357);
  not g29915 (n_14358, n15776);
  and g29916 (n15816, n_14358, n15814);
  and g29917 (n15817, n15647, n15706);
  not g29918 (n_14359, n15647);
  not g29919 (n_14360, n15706);
  and g29920 (n15818, n_14359, n_14360);
  not g29921 (n_14361, n15817);
  not g29922 (n_14362, n15818);
  and g29923 (n15819, n_14361, n_14362);
  and g29924 (n15820, n_14263, n_14270);
  not g29925 (n_14363, n15819);
  and g29926 (n15821, n_14363, n15820);
  not g29927 (n_14364, n15820);
  and g29928 (n15822, n15819, n_14364);
  not g29929 (n_14365, n15821);
  not g29930 (n_14366, n15822);
  and g29931 (n15823, n_14365, n_14366);
  and g29932 (n15824, n_14244, n_14250);
  not g29933 (n_14367, n15823);
  and g29934 (n15825, n_14367, n15824);
  not g29935 (n_14368, n15824);
  and g29936 (n15826, n15823, n_14368);
  not g29937 (n_14369, n15825);
  not g29938 (n_14370, n15826);
  and g29939 (n15827, n_14369, n_14370);
  and g29940 (n15828, \a[40] , \a[51] );
  and g29941 (n15829, \a[41] , \a[50] );
  not g29942 (n_14371, n15828);
  not g29943 (n_14372, n15829);
  and g29944 (n15830, n_14371, n_14372);
  and g29945 (n15831, n5413, n6564);
  not g29946 (n_14373, n15831);
  not g29949 (n_14374, n15830);
  not g29951 (n_14375, n15834);
  and g29952 (n15835, n_14373, n_14375);
  and g29953 (n15836, n_14374, n15835);
  and g29954 (n15837, \a[63] , n_14375);
  and g29955 (n15838, \a[28] , n15837);
  not g29956 (n_14376, n15836);
  not g29957 (n_14377, n15838);
  and g29958 (n15839, n_14376, n_14377);
  and g29959 (n15840, \a[43] , \a[48] );
  and g29960 (n15841, \a[44] , \a[47] );
  not g29961 (n_14378, n15840);
  not g29962 (n_14379, n15841);
  and g29963 (n15842, n_14378, n_14379);
  and g29964 (n15843, n5296, n6252);
  not g29965 (n_14380, n15843);
  not g29968 (n_14381, n15842);
  not g29970 (n_14382, n15846);
  and g29971 (n15847, \a[56] , n_14382);
  and g29972 (n15848, \a[35] , n15847);
  and g29973 (n15849, n_14380, n_14382);
  and g29974 (n15850, n_14381, n15849);
  not g29975 (n_14383, n15848);
  not g29976 (n_14384, n15850);
  and g29977 (n15851, n_14383, n_14384);
  not g29978 (n_14385, n15839);
  not g29979 (n_14386, n15851);
  and g29980 (n15852, n_14385, n_14386);
  not g29981 (n_14387, n15852);
  and g29982 (n15853, n_14385, n_14387);
  and g29983 (n15854, n_14386, n_14387);
  not g29984 (n_14388, n15853);
  not g29985 (n_14389, n15854);
  and g29986 (n15855, n_14388, n_14389);
  and g29987 (n15856, \a[46] , \a[62] );
  and g29988 (n15857, \a[29] , n15856);
  not g29989 (n_14390, n15857);
  and g29990 (n15858, n5560, n_14390);
  not g29991 (n_14391, n15858);
  and g29992 (n15859, n5560, n_14391);
  and g29993 (n15860, n_14390, n_14391);
  and g29994 (n15861, \a[29] , \a[62] );
  not g29995 (n_14392, \a[46] );
  not g29996 (n_14393, n15861);
  and g29997 (n15862, n_14392, n_14393);
  not g29998 (n_14394, n15862);
  and g29999 (n15863, n15860, n_14394);
  not g30000 (n_14395, n15859);
  not g30001 (n_14396, n15863);
  and g30002 (n15864, n_14395, n_14396);
  not g30003 (n_14397, n15855);
  not g30004 (n_14398, n15864);
  and g30005 (n15865, n_14397, n_14398);
  not g30006 (n_14399, n15865);
  and g30007 (n15866, n_14397, n_14399);
  and g30008 (n15867, n_14398, n_14399);
  not g30009 (n_14400, n15866);
  not g30010 (n_14401, n15867);
  and g30011 (n15868, n_14400, n_14401);
  not g30012 (n_14402, n15827);
  and g30013 (n15869, n_14402, n15868);
  not g30014 (n_14403, n15868);
  and g30015 (n15870, n15827, n_14403);
  not g30016 (n_14404, n15869);
  not g30017 (n_14405, n15870);
  and g30018 (n15871, n_14404, n_14405);
  and g30019 (n15872, n_14162, n_14167);
  not g30020 (n_14406, n15872);
  and g30021 (n15873, n15871, n_14406);
  not g30022 (n_14407, n15871);
  and g30023 (n15874, n_14407, n15872);
  not g30024 (n_14408, n15873);
  not g30025 (n_14409, n15874);
  and g30026 (n15875, n_14408, n_14409);
  not g30027 (n_14410, n15816);
  and g30028 (n15876, n_14410, n15875);
  not g30029 (n_14411, n15815);
  and g30030 (n15877, n_14411, n15876);
  not g30031 (n_14412, n15877);
  and g30032 (n15878, n15875, n_14412);
  and g30033 (n15879, n_14410, n_14412);
  and g30034 (n15880, n_14411, n15879);
  not g30035 (n_14413, n15878);
  not g30036 (n_14414, n15880);
  and g30037 (n15881, n_14413, n_14414);
  and g30038 (n15882, n_14229, n_14290);
  and g30039 (n15883, n_14280, n_14285);
  and g30040 (n15884, n_14183, n_14228);
  and g30041 (n15885, \a[30] , \a[61] );
  not g30042 (n_14415, n15663);
  and g30043 (n15886, n_14415, n15885);
  not g30044 (n_14416, n15885);
  and g30045 (n15887, n15663, n_14416);
  not g30046 (n_14417, n15886);
  not g30047 (n_14418, n15887);
  and g30048 (n15888, n_14417, n_14418);
  not g30049 (n_14419, n15888);
  and g30050 (n15889, n15635, n_14419);
  not g30051 (n_14420, n15635);
  and g30052 (n15890, n_14420, n15888);
  not g30053 (n_14421, n15889);
  not g30054 (n_14422, n15890);
  and g30055 (n15891, n_14421, n_14422);
  and g30056 (n15892, n_14273, n_14278);
  and g30057 (n15893, n_14206, n_14221);
  and g30058 (n15894, n15892, n15893);
  not g30059 (n_14423, n15892);
  not g30060 (n_14424, n15893);
  and g30061 (n15895, n_14423, n_14424);
  not g30062 (n_14425, n15894);
  not g30063 (n_14426, n15895);
  and g30064 (n15896, n_14425, n_14426);
  and g30065 (n15897, n15891, n15896);
  not g30066 (n_14427, n15891);
  not g30067 (n_14428, n15896);
  and g30068 (n15898, n_14427, n_14428);
  not g30069 (n_14429, n15897);
  not g30070 (n_14430, n15898);
  and g30071 (n15899, n_14429, n_14430);
  not g30072 (n_14431, n15884);
  and g30073 (n15900, n_14431, n15899);
  not g30074 (n_14432, n15900);
  and g30075 (n15901, n_14431, n_14432);
  and g30076 (n15902, n15899, n_14432);
  not g30077 (n_14433, n15901);
  not g30078 (n_14434, n15902);
  and g30079 (n15903, n_14433, n_14434);
  not g30080 (n_14435, n15883);
  not g30081 (n_14436, n15903);
  and g30082 (n15904, n_14435, n_14436);
  not g30083 (n_14437, n15904);
  and g30084 (n15905, n_14435, n_14437);
  and g30085 (n15906, n_14436, n_14437);
  not g30086 (n_14438, n15905);
  not g30087 (n_14439, n15906);
  and g30088 (n15907, n_14438, n_14439);
  not g30089 (n_14440, n15882);
  not g30090 (n_14441, n15907);
  and g30091 (n15908, n_14440, n_14441);
  not g30092 (n_14442, n15908);
  and g30093 (n15909, n_14440, n_14442);
  and g30094 (n15910, n_14441, n_14442);
  not g30095 (n_14443, n15909);
  not g30096 (n_14444, n15910);
  and g30097 (n15911, n_14443, n_14444);
  not g30098 (n_14445, n15881);
  and g30099 (n15912, n_14445, n15911);
  not g30100 (n_14446, n15911);
  and g30101 (n15913, n15881, n_14446);
  not g30102 (n_14447, n15912);
  not g30103 (n_14448, n15913);
  and g30104 (n15914, n_14447, n_14448);
  not g30105 (n_14449, n15757);
  not g30106 (n_14450, n15914);
  and g30107 (n15915, n_14449, n_14450);
  and g30108 (n15916, n15757, n15914);
  not g30109 (n_14451, n15915);
  not g30110 (n_14452, n15916);
  and g30111 (n15917, n_14451, n_14452);
  not g30112 (n_14453, n15756);
  not g30113 (n_14454, n15917);
  and g30114 (n15918, n_14453, n_14454);
  and g30115 (n15919, n15756, n15917);
  or g30116 (\asquared[92] , n15918, n15919);
  and g30117 (n15921, n_14453, n_14452);
  not g30118 (n_14455, n15921);
  and g30119 (n15922, n_14451, n_14455);
  and g30120 (n15923, n_14432, n_14437);
  and g30121 (n15924, n_14354, n_14411);
  and g30122 (n15925, n_14426, n_14429);
  and g30123 (n15926, n2865, n9721);
  not g30124 (n_14456, n15926);
  and g30125 (n15927, \a[61] , n_14456);
  and g30126 (n15928, \a[31] , n15927);
  and g30127 (n15929, \a[62] , n_14456);
  and g30128 (n15930, \a[30] , n15929);
  not g30129 (n_14457, n15928);
  not g30130 (n_14458, n15930);
  and g30131 (n15931, n_14457, n_14458);
  not g30132 (n_14459, n15860);
  not g30133 (n_14460, n15931);
  and g30134 (n15932, n_14459, n_14460);
  not g30135 (n_14461, n15932);
  and g30136 (n15933, n_14459, n_14461);
  and g30137 (n15934, n_14460, n_14461);
  not g30138 (n_14462, n15933);
  not g30139 (n_14463, n15934);
  and g30140 (n15935, n_14462, n_14463);
  and g30141 (n15936, n5413, n6968);
  and g30142 (n15937, n3984, n7232);
  and g30143 (n15938, n4171, n7433);
  not g30144 (n_14464, n15937);
  not g30145 (n_14465, n15938);
  and g30146 (n15939, n_14464, n_14465);
  not g30147 (n_14466, n15936);
  not g30148 (n_14467, n15939);
  and g30149 (n15940, n_14466, n_14467);
  not g30150 (n_14468, n15940);
  and g30151 (n15941, \a[53] , n_14468);
  and g30152 (n15942, \a[39] , n15941);
  and g30153 (n15943, \a[40] , \a[52] );
  and g30154 (n15944, \a[41] , \a[51] );
  not g30155 (n_14469, n15943);
  not g30156 (n_14470, n15944);
  and g30157 (n15945, n_14469, n_14470);
  and g30158 (n15946, n_14466, n_14468);
  not g30159 (n_14471, n15945);
  and g30160 (n15947, n_14471, n15946);
  not g30161 (n_14472, n15942);
  not g30162 (n_14473, n15947);
  and g30163 (n15948, n_14472, n_14473);
  not g30164 (n_14474, n15935);
  not g30165 (n_14475, n15948);
  and g30166 (n15949, n_14474, n_14475);
  not g30167 (n_14476, n15949);
  and g30168 (n15950, n_14474, n_14476);
  and g30169 (n15951, n_14475, n_14476);
  not g30170 (n_14477, n15950);
  not g30171 (n_14478, n15951);
  and g30172 (n15952, n_14477, n_14478);
  and g30173 (n15953, n_14417, n_14422);
  and g30174 (n15954, n15952, n15953);
  not g30175 (n_14479, n15952);
  not g30176 (n_14480, n15953);
  and g30177 (n15955, n_14479, n_14480);
  not g30178 (n_14481, n15954);
  not g30179 (n_14482, n15955);
  and g30180 (n15956, n_14481, n_14482);
  and g30181 (n15957, \a[42] , \a[50] );
  and g30182 (n15958, \a[34] , n15957);
  and g30183 (n15959, \a[58] , n15958);
  and g30184 (n15960, n3319, n8436);
  not g30185 (n_14483, n15959);
  not g30186 (n_14484, n15960);
  and g30187 (n15961, n_14483, n_14484);
  and g30188 (n15962, \a[35] , \a[57] );
  and g30189 (n15963, n15957, n15962);
  not g30190 (n_14485, n15961);
  not g30191 (n_14486, n15963);
  and g30192 (n15964, n_14485, n_14486);
  not g30193 (n_14487, n15964);
  and g30194 (n15965, n_14486, n_14487);
  not g30195 (n_14488, n15957);
  not g30196 (n_14489, n15962);
  and g30197 (n15966, n_14488, n_14489);
  not g30198 (n_14490, n15966);
  and g30199 (n15967, n15965, n_14490);
  and g30200 (n15968, \a[58] , n_14487);
  and g30201 (n15969, \a[34] , n15968);
  not g30202 (n_14491, n15967);
  not g30203 (n_14492, n15969);
  and g30204 (n15970, n_14491, n_14492);
  and g30205 (n15971, n5713, n6252);
  and g30206 (n15972, n4811, n6254);
  and g30207 (n15973, n5296, n6256);
  not g30208 (n_14493, n15972);
  not g30209 (n_14494, n15973);
  and g30210 (n15974, n_14493, n_14494);
  not g30211 (n_14495, n15971);
  not g30212 (n_14496, n15974);
  and g30213 (n15975, n_14495, n_14496);
  not g30214 (n_14497, n15975);
  and g30215 (n15976, \a[49] , n_14497);
  and g30216 (n15977, \a[43] , n15976);
  and g30217 (n15978, n_14495, n_14497);
  and g30218 (n15979, \a[44] , \a[48] );
  not g30219 (n_14498, n5250);
  not g30220 (n_14499, n15979);
  and g30221 (n15980, n_14498, n_14499);
  not g30222 (n_14500, n15980);
  and g30223 (n15981, n15978, n_14500);
  not g30224 (n_14501, n15977);
  not g30225 (n_14502, n15981);
  and g30226 (n15982, n_14501, n_14502);
  not g30227 (n_14503, n15970);
  not g30228 (n_14504, n15982);
  and g30229 (n15983, n_14503, n_14504);
  not g30230 (n_14505, n15983);
  and g30231 (n15984, n_14503, n_14505);
  and g30232 (n15985, n_14504, n_14505);
  not g30233 (n_14506, n15984);
  not g30234 (n_14507, n15985);
  and g30235 (n15986, n_14506, n_14507);
  and g30236 (n15987, \a[36] , \a[56] );
  and g30237 (n15988, \a[33] , \a[59] );
  not g30238 (n_14508, n13656);
  not g30239 (n_14509, n15988);
  and g30240 (n15989, n_14508, n_14509);
  and g30241 (n15990, n13656, n15988);
  not g30242 (n_14510, n15990);
  and g30243 (n15991, n15987, n_14510);
  not g30244 (n_14511, n15989);
  and g30245 (n15992, n_14511, n15991);
  not g30246 (n_14512, n15992);
  and g30247 (n15993, n15987, n_14512);
  and g30248 (n15994, n_14510, n_14512);
  and g30249 (n15995, n_14511, n15994);
  not g30250 (n_14513, n15993);
  not g30251 (n_14514, n15995);
  and g30252 (n15996, n_14513, n_14514);
  not g30253 (n_14515, n15986);
  not g30254 (n_14516, n15996);
  and g30255 (n15997, n_14515, n_14516);
  not g30256 (n_14517, n15997);
  and g30257 (n15998, n_14515, n_14517);
  and g30258 (n15999, n_14516, n_14517);
  not g30259 (n_14518, n15998);
  not g30260 (n_14519, n15999);
  and g30261 (n16000, n_14518, n_14519);
  not g30262 (n_14520, n15956);
  and g30263 (n16001, n_14520, n16000);
  not g30264 (n_14521, n16000);
  and g30265 (n16002, n15956, n_14521);
  not g30266 (n_14522, n16001);
  not g30267 (n_14523, n16002);
  and g30268 (n16003, n_14522, n_14523);
  not g30269 (n_14524, n15925);
  and g30270 (n16004, n_14524, n16003);
  not g30271 (n_14525, n16003);
  and g30272 (n16005, n15925, n_14525);
  not g30273 (n_14526, n16004);
  not g30274 (n_14527, n16005);
  and g30275 (n16006, n_14526, n_14527);
  not g30276 (n_14528, n15924);
  and g30277 (n16007, n_14528, n16006);
  not g30278 (n_14529, n16006);
  and g30279 (n16008, n15924, n_14529);
  not g30280 (n_14530, n16007);
  not g30281 (n_14531, n16008);
  and g30282 (n16009, n_14530, n_14531);
  not g30283 (n_14532, n15923);
  and g30284 (n16010, n_14532, n16009);
  not g30285 (n_14533, n16009);
  and g30286 (n16011, n15923, n_14533);
  not g30287 (n_14534, n16010);
  not g30288 (n_14535, n16011);
  and g30289 (n16012, n_14534, n_14535);
  and g30290 (n16013, n_14408, n_14412);
  and g30291 (n16014, n_14344, n_14349);
  and g30292 (n16015, n_14362, n_14366);
  and g30293 (n16016, n16014, n16015);
  not g30294 (n_14536, n16014);
  not g30295 (n_14537, n16015);
  and g30296 (n16017, n_14536, n_14537);
  not g30297 (n_14538, n16016);
  not g30298 (n_14539, n16017);
  and g30299 (n16018, n_14538, n_14539);
  and g30300 (n16019, n_14387, n_14399);
  not g30301 (n_14540, n16018);
  and g30302 (n16020, n_14540, n16019);
  not g30303 (n_14541, n16019);
  and g30304 (n16021, n16018, n_14541);
  not g30305 (n_14542, n16020);
  not g30306 (n_14543, n16021);
  and g30307 (n16022, n_14542, n_14543);
  and g30308 (n16023, n_14370, n_14405);
  and g30309 (n16024, n_14315, n_14321);
  and g30310 (n16025, n15783, n15797);
  not g30311 (n_14544, n15783);
  not g30312 (n_14545, n15797);
  and g30313 (n16026, n_14544, n_14545);
  not g30314 (n_14546, n16025);
  not g30315 (n_14547, n16026);
  and g30316 (n16027, n_14546, n_14547);
  not g30317 (n_14548, n16027);
  and g30318 (n16028, n15835, n_14548);
  not g30319 (n_14549, n15835);
  and g30320 (n16029, n_14549, n16027);
  not g30321 (n_14550, n16028);
  not g30322 (n_14551, n16029);
  and g30323 (n16030, n_14550, n_14551);
  and g30324 (n16031, n15766, n15849);
  not g30325 (n_14552, n15766);
  not g30326 (n_14553, n15849);
  and g30327 (n16032, n_14552, n_14553);
  not g30328 (n_14554, n16031);
  not g30329 (n_14555, n16032);
  and g30330 (n16033, n_14554, n_14555);
  and g30331 (n16034, n4565, n7701);
  and g30332 (n16035, \a[37] , \a[55] );
  and g30333 (n16036, \a[38] , \a[54] );
  not g30334 (n_14556, n16035);
  not g30335 (n_14557, n16036);
  and g30336 (n16037, n_14556, n_14557);
  not g30337 (n_14558, n16034);
  not g30338 (n_14559, n16037);
  not g30342 (n_14560, n16040);
  and g30343 (n16041, \a[60] , n_14560);
  and g30344 (n16042, \a[32] , n16041);
  and g30345 (n16043, n_14558, n_14560);
  and g30346 (n16044, n_14559, n16043);
  not g30347 (n_14561, n16042);
  not g30348 (n_14562, n16044);
  and g30349 (n16045, n_14561, n_14562);
  not g30350 (n_14563, n16045);
  and g30351 (n16046, n16033, n_14563);
  not g30352 (n_14564, n16046);
  and g30353 (n16047, n16033, n_14564);
  and g30354 (n16048, n_14563, n_14564);
  not g30355 (n_14565, n16047);
  not g30356 (n_14566, n16048);
  and g30357 (n16049, n_14565, n_14566);
  not g30358 (n_14567, n16030);
  and g30359 (n16050, n_14567, n16049);
  not g30360 (n_14568, n16049);
  and g30361 (n16051, n16030, n_14568);
  not g30362 (n_14569, n16050);
  not g30363 (n_14570, n16051);
  and g30364 (n16052, n_14569, n_14570);
  not g30365 (n_14571, n16024);
  and g30366 (n16053, n_14571, n16052);
  not g30367 (n_14572, n16052);
  and g30368 (n16054, n16024, n_14572);
  not g30369 (n_14573, n16053);
  not g30370 (n_14574, n16054);
  and g30371 (n16055, n_14573, n_14574);
  not g30372 (n_14575, n16023);
  and g30373 (n16056, n_14575, n16055);
  not g30374 (n_14576, n16055);
  and g30375 (n16057, n16023, n_14576);
  not g30376 (n_14577, n16056);
  not g30377 (n_14578, n16057);
  and g30378 (n16058, n_14577, n_14578);
  and g30379 (n16059, n16022, n16058);
  not g30380 (n_14579, n16022);
  not g30381 (n_14580, n16058);
  and g30382 (n16060, n_14579, n_14580);
  not g30383 (n_14581, n16059);
  not g30384 (n_14582, n16060);
  and g30385 (n16061, n_14581, n_14582);
  not g30386 (n_14583, n16013);
  and g30387 (n16062, n_14583, n16061);
  not g30388 (n_14584, n16061);
  and g30389 (n16063, n16013, n_14584);
  not g30390 (n_14585, n16062);
  not g30391 (n_14586, n16063);
  and g30392 (n16064, n_14585, n_14586);
  and g30393 (n16065, n16012, n16064);
  not g30394 (n_14587, n16012);
  not g30395 (n_14588, n16064);
  and g30396 (n16066, n_14587, n_14588);
  not g30397 (n_14589, n16065);
  not g30398 (n_14590, n16066);
  and g30399 (n16067, n_14589, n_14590);
  and g30400 (n16068, n_14445, n_14446);
  not g30401 (n_14591, n16068);
  and g30402 (n16069, n_14442, n_14591);
  not g30403 (n_14592, n16067);
  and g30404 (n16070, n_14592, n16069);
  not g30405 (n_14593, n16069);
  and g30406 (n16071, n16067, n_14593);
  not g30407 (n_14594, n16070);
  not g30408 (n_14595, n16071);
  and g30409 (n16072, n_14594, n_14595);
  not g30410 (n_14596, n16072);
  and g30411 (n16073, n15922, n_14596);
  not g30412 (n_14597, n15922);
  and g30413 (n16074, n_14597, n_14594);
  and g30414 (n16075, n_14595, n16074);
  not g30415 (n_14598, n16073);
  not g30416 (n_14599, n16075);
  and g30417 (\asquared[93] , n_14598, n_14599);
  not g30418 (n_14600, n16074);
  and g30419 (n16077, n_14595, n_14600);
  and g30420 (n16078, n_14585, n_14589);
  and g30421 (n16079, n_14530, n_14534);
  and g30422 (n16080, n_14555, n_14564);
  and g30423 (n16081, n_14547, n_14551);
  and g30424 (n16082, n16080, n16081);
  not g30425 (n_14601, n16080);
  not g30426 (n_14602, n16081);
  and g30427 (n16083, n_14601, n_14602);
  not g30428 (n_14603, n16082);
  not g30429 (n_14604, n16083);
  and g30430 (n16084, n_14603, n_14604);
  and g30431 (n16085, n_14505, n_14517);
  not g30432 (n_14605, n16084);
  and g30433 (n16086, n_14605, n16085);
  not g30434 (n_14606, n16085);
  and g30435 (n16087, n16084, n_14606);
  not g30436 (n_14607, n16086);
  not g30437 (n_14608, n16087);
  and g30438 (n16088, n_14607, n_14608);
  and g30439 (n16089, n_14570, n_14573);
  not g30440 (n_14609, n16089);
  and g30441 (n16090, n16088, n_14609);
  not g30442 (n_14610, n16088);
  and g30443 (n16091, n_14610, n16089);
  not g30444 (n_14611, n16090);
  not g30445 (n_14612, n16091);
  and g30446 (n16092, n_14611, n_14612);
  and g30447 (n16093, n_14476, n_14482);
  and g30448 (n16094, n15965, n15978);
  not g30449 (n_14613, n15965);
  not g30450 (n_14614, n15978);
  and g30451 (n16095, n_14613, n_14614);
  not g30452 (n_14615, n16094);
  not g30453 (n_14616, n16095);
  and g30454 (n16096, n_14615, n_14616);
  not g30455 (n_14617, n16096);
  and g30456 (n16097, n15946, n_14617);
  not g30457 (n_14618, n15946);
  and g30458 (n16098, n_14618, n16096);
  not g30459 (n_14619, n16097);
  not g30460 (n_14620, n16098);
  and g30461 (n16099, n_14619, n_14620);
  and g30462 (n16100, n15994, n16043);
  not g30463 (n_14621, n15994);
  not g30464 (n_14622, n16043);
  and g30465 (n16101, n_14621, n_14622);
  not g30466 (n_14623, n16100);
  not g30467 (n_14624, n16101);
  and g30468 (n16102, n_14623, n_14624);
  and g30469 (n16103, n_14456, n_14461);
  not g30470 (n_14625, n16102);
  and g30471 (n16104, n_14625, n16103);
  not g30472 (n_14626, n16103);
  and g30473 (n16105, n16102, n_14626);
  not g30474 (n_14627, n16104);
  not g30475 (n_14628, n16105);
  and g30476 (n16106, n_14627, n_14628);
  and g30477 (n16107, n16099, n16106);
  not g30478 (n_14629, n16099);
  not g30479 (n_14630, n16106);
  and g30480 (n16108, n_14629, n_14630);
  not g30481 (n_14631, n16107);
  not g30482 (n_14632, n16108);
  and g30483 (n16109, n_14631, n_14632);
  not g30484 (n_14633, n16093);
  and g30485 (n16110, n_14633, n16109);
  not g30486 (n_14634, n16109);
  and g30487 (n16111, n16093, n_14634);
  not g30488 (n_14635, n16110);
  not g30489 (n_14636, n16111);
  and g30490 (n16112, n_14635, n_14636);
  and g30491 (n16113, n16092, n16112);
  not g30492 (n_14637, n16092);
  not g30493 (n_14638, n16112);
  and g30494 (n16114, n_14637, n_14638);
  not g30495 (n_14639, n16113);
  not g30496 (n_14640, n16114);
  and g30497 (n16115, n_14639, n_14640);
  not g30498 (n_14641, n16115);
  and g30499 (n16116, n16079, n_14641);
  not g30500 (n_14642, n16079);
  and g30501 (n16117, n_14642, n16115);
  not g30502 (n_14643, n16116);
  not g30503 (n_14644, n16117);
  and g30504 (n16118, n_14643, n_14644);
  and g30505 (n16119, n_14577, n_14581);
  and g30506 (n16120, n_14523, n_14526);
  and g30507 (n16121, n_14539, n_14543);
  and g30508 (n16122, n3143, n9512);
  and g30509 (n16123, n9475, n11634);
  and g30510 (n16124, n2488, n9909);
  not g30511 (n_14645, n16123);
  not g30512 (n_14646, n16124);
  and g30513 (n16125, n_14645, n_14646);
  not g30514 (n_14647, n16122);
  not g30515 (n_14648, n16125);
  and g30516 (n16126, n_14647, n_14648);
  not g30517 (n_14649, n16126);
  and g30518 (n16127, n_14647, n_14649);
  and g30519 (n16128, \a[32] , \a[61] );
  and g30520 (n16129, \a[33] , \a[60] );
  not g30521 (n_14650, n16128);
  not g30522 (n_14651, n16129);
  and g30523 (n16130, n_14650, n_14651);
  not g30524 (n_14652, n16130);
  and g30525 (n16131, n16127, n_14652);
  and g30526 (n16132, \a[63] , n_14649);
  and g30527 (n16133, \a[30] , n16132);
  not g30528 (n_14653, n16131);
  not g30529 (n_14654, n16133);
  and g30530 (n16134, n_14653, n_14654);
  and g30531 (n16135, n8936, n13730);
  and g30532 (n16136, n3828, n8436);
  and g30533 (n16137, \a[39] , \a[54] );
  and g30534 (n16138, n15203, n16137);
  not g30535 (n_14655, n16136);
  not g30536 (n_14656, n16138);
  and g30537 (n16139, n_14655, n_14656);
  not g30538 (n_14657, n16135);
  not g30539 (n_14658, n16139);
  and g30540 (n16140, n_14657, n_14658);
  not g30541 (n_14659, n16140);
  and g30542 (n16141, n15203, n_14659);
  and g30543 (n16142, n_14657, n_14659);
  and g30544 (n16143, \a[36] , \a[57] );
  not g30545 (n_14660, n16137);
  not g30546 (n_14661, n16143);
  and g30547 (n16144, n_14660, n_14661);
  not g30548 (n_14662, n16144);
  and g30549 (n16145, n16142, n_14662);
  not g30550 (n_14663, n16141);
  not g30551 (n_14664, n16145);
  and g30552 (n16146, n_14663, n_14664);
  not g30553 (n_14665, n16134);
  not g30554 (n_14666, n16146);
  and g30555 (n16147, n_14665, n_14666);
  not g30556 (n_14667, n16147);
  and g30557 (n16148, n_14665, n_14667);
  and g30558 (n16149, n_14666, n_14667);
  not g30559 (n_14668, n16148);
  not g30560 (n_14669, n16149);
  and g30561 (n16150, n_14668, n_14669);
  and g30562 (n16151, \a[40] , \a[53] );
  and g30563 (n16152, \a[41] , \a[52] );
  not g30564 (n_14670, n16151);
  not g30565 (n_14671, n16152);
  and g30566 (n16153, n_14670, n_14671);
  and g30567 (n16154, n5413, n7433);
  not g30568 (n_14672, n16154);
  and g30569 (n16155, n15188, n_14672);
  not g30570 (n_14673, n16153);
  and g30571 (n16156, n_14673, n16155);
  not g30572 (n_14674, n16156);
  and g30573 (n16157, n15188, n_14674);
  and g30574 (n16158, n_14672, n_14674);
  and g30575 (n16159, n_14673, n16158);
  not g30576 (n_14675, n16157);
  not g30577 (n_14676, n16159);
  and g30578 (n16160, n_14675, n_14676);
  not g30579 (n_14677, n16150);
  not g30580 (n_14678, n16160);
  and g30581 (n16161, n_14677, n_14678);
  not g30582 (n_14679, n16161);
  and g30583 (n16162, n_14677, n_14679);
  and g30584 (n16163, n_14678, n_14679);
  not g30585 (n_14680, n16162);
  not g30586 (n_14681, n16163);
  and g30587 (n16164, n_14680, n_14681);
  and g30588 (n16165, \a[38] , \a[55] );
  not g30589 (n_14682, n8155);
  not g30590 (n_14683, n16165);
  and g30591 (n16166, n_14682, n_14683);
  and g30592 (n16167, \a[45] , \a[55] );
  and g30593 (n16168, n6942, n16167);
  and g30594 (n16169, n6146, n9666);
  and g30595 (n16170, n4565, n9161);
  not g30596 (n_14684, n16169);
  not g30597 (n_14685, n16170);
  and g30598 (n16171, n_14684, n_14685);
  not g30599 (n_14686, n16168);
  not g30600 (n_14687, n16171);
  and g30601 (n16172, n_14686, n_14687);
  not g30602 (n_14688, n16172);
  and g30603 (n16173, n_14686, n_14688);
  not g30604 (n_14689, n16166);
  and g30605 (n16174, n_14689, n16173);
  and g30606 (n16175, \a[56] , n_14688);
  and g30607 (n16176, \a[37] , n16175);
  not g30608 (n_14690, n16174);
  not g30609 (n_14691, n16176);
  and g30610 (n16177, n_14690, n_14691);
  and g30611 (n16178, n5296, n6325);
  and g30612 (n16179, n4639, n9934);
  and g30613 (n16180, n5018, n6564);
  not g30614 (n_14692, n16179);
  not g30615 (n_14693, n16180);
  and g30616 (n16181, n_14692, n_14693);
  not g30617 (n_14694, n16178);
  not g30618 (n_14695, n16181);
  and g30619 (n16182, n_14694, n_14695);
  not g30620 (n_14696, n16182);
  and g30621 (n16183, \a[51] , n_14696);
  and g30622 (n16184, \a[42] , n16183);
  and g30623 (n16185, n_14694, n_14696);
  and g30624 (n16186, \a[43] , \a[50] );
  not g30625 (n_14697, n8252);
  not g30626 (n_14698, n16186);
  and g30627 (n16187, n_14697, n_14698);
  not g30628 (n_14699, n16187);
  and g30629 (n16188, n16185, n_14699);
  not g30630 (n_14700, n16184);
  not g30631 (n_14701, n16188);
  and g30632 (n16189, n_14700, n_14701);
  not g30633 (n_14702, n16177);
  not g30634 (n_14703, n16189);
  and g30635 (n16190, n_14702, n_14703);
  not g30636 (n_14704, n16190);
  and g30637 (n16191, n_14702, n_14704);
  and g30638 (n16192, n_14703, n_14704);
  not g30639 (n_14705, n16191);
  not g30640 (n_14706, n16192);
  and g30641 (n16193, n_14705, n_14706);
  and g30642 (n16194, \a[47] , \a[62] );
  and g30643 (n16195, \a[31] , n16194);
  not g30644 (n_14707, n16195);
  and g30645 (n16196, n5666, n_14707);
  not g30646 (n_14708, n16196);
  and g30647 (n16197, n5666, n_14708);
  and g30648 (n16198, n_14707, n_14708);
  and g30649 (n16199, \a[31] , \a[62] );
  not g30650 (n_14709, \a[47] );
  not g30651 (n_14710, n16199);
  and g30652 (n16200, n_14709, n_14710);
  not g30653 (n_14711, n16200);
  and g30654 (n16201, n16198, n_14711);
  not g30655 (n_14712, n16197);
  not g30656 (n_14713, n16201);
  and g30657 (n16202, n_14712, n_14713);
  not g30658 (n_14714, n16193);
  not g30659 (n_14715, n16202);
  and g30660 (n16203, n_14714, n_14715);
  not g30661 (n_14716, n16203);
  and g30662 (n16204, n_14714, n_14716);
  and g30663 (n16205, n_14715, n_14716);
  not g30664 (n_14717, n16204);
  not g30665 (n_14718, n16205);
  and g30666 (n16206, n_14717, n_14718);
  and g30667 (n16207, n16164, n16206);
  not g30668 (n_14719, n16164);
  not g30669 (n_14720, n16206);
  and g30670 (n16208, n_14719, n_14720);
  not g30671 (n_14721, n16207);
  not g30672 (n_14722, n16208);
  and g30673 (n16209, n_14721, n_14722);
  not g30674 (n_14723, n16121);
  and g30675 (n16210, n_14723, n16209);
  not g30676 (n_14724, n16209);
  and g30677 (n16211, n16121, n_14724);
  not g30678 (n_14725, n16210);
  not g30679 (n_14726, n16211);
  and g30680 (n16212, n_14725, n_14726);
  not g30681 (n_14727, n16120);
  and g30682 (n16213, n_14727, n16212);
  not g30683 (n_14728, n16212);
  and g30684 (n16214, n16120, n_14728);
  not g30685 (n_14729, n16213);
  not g30686 (n_14730, n16214);
  and g30687 (n16215, n_14729, n_14730);
  not g30688 (n_14731, n16215);
  and g30689 (n16216, n16119, n_14731);
  not g30690 (n_14732, n16119);
  and g30691 (n16217, n_14732, n16215);
  not g30692 (n_14733, n16216);
  not g30693 (n_14734, n16217);
  and g30694 (n16218, n_14733, n_14734);
  and g30695 (n16219, n16118, n16218);
  not g30696 (n_14735, n16118);
  not g30697 (n_14736, n16218);
  and g30698 (n16220, n_14735, n_14736);
  not g30699 (n_14737, n16219);
  not g30700 (n_14738, n16220);
  and g30701 (n16221, n_14737, n_14738);
  not g30702 (n_14739, n16078);
  and g30703 (n16222, n_14739, n16221);
  not g30704 (n_14740, n16221);
  and g30705 (n16223, n16078, n_14740);
  not g30706 (n_14741, n16222);
  not g30707 (n_14742, n16223);
  and g30708 (n16224, n_14741, n_14742);
  not g30709 (n_14743, n16077);
  not g30710 (n_14744, n16224);
  and g30711 (n16225, n_14743, n_14744);
  and g30712 (n16226, n16077, n16224);
  or g30713 (\asquared[94] , n16225, n16226);
  and g30714 (n16228, n_14729, n_14734);
  and g30715 (n16229, n_14722, n_14725);
  and g30716 (n16230, n_14624, n_14628);
  and g30717 (n16231, n_14616, n_14620);
  and g30718 (n16232, n16230, n16231);
  not g30719 (n_14745, n16230);
  not g30720 (n_14746, n16231);
  and g30721 (n16233, n_14745, n_14746);
  not g30722 (n_14747, n16232);
  not g30723 (n_14748, n16233);
  and g30724 (n16234, n_14747, n_14748);
  and g30725 (n16235, n_14667, n_14679);
  not g30726 (n_14749, n16234);
  and g30727 (n16236, n_14749, n16235);
  not g30728 (n_14750, n16235);
  and g30729 (n16237, n16234, n_14750);
  not g30730 (n_14751, n16236);
  not g30731 (n_14752, n16237);
  and g30732 (n16238, n_14751, n_14752);
  and g30733 (n16239, n_14631, n_14635);
  not g30734 (n_14753, n16239);
  and g30735 (n16240, n16238, n_14753);
  not g30736 (n_14754, n16238);
  and g30737 (n16241, n_14754, n16239);
  not g30738 (n_14755, n16240);
  not g30739 (n_14756, n16241);
  and g30740 (n16242, n_14755, n_14756);
  not g30741 (n_14757, n16229);
  and g30742 (n16243, n_14757, n16242);
  not g30743 (n_14758, n16242);
  and g30744 (n16244, n16229, n_14758);
  not g30745 (n_14759, n16243);
  not g30746 (n_14760, n16244);
  and g30747 (n16245, n_14759, n_14760);
  not g30748 (n_14761, n16245);
  and g30749 (n16246, n16228, n_14761);
  not g30750 (n_14762, n16228);
  and g30751 (n16247, n_14762, n16245);
  not g30752 (n_14763, n16246);
  not g30753 (n_14764, n16247);
  and g30754 (n16248, n_14763, n_14764);
  and g30755 (n16249, \a[43] , \a[51] );
  not g30756 (n_14765, n8254);
  not g30757 (n_14766, n16249);
  and g30758 (n16250, n_14765, n_14766);
  and g30759 (n16251, n5296, n6564);
  not g30760 (n_14767, n16251);
  not g30763 (n_14768, n16250);
  not g30765 (n_14769, n16254);
  and g30766 (n16255, n_14767, n_14769);
  and g30767 (n16256, n_14768, n16255);
  and g30768 (n16257, \a[58] , n_14769);
  and g30769 (n16258, \a[36] , n16257);
  not g30770 (n_14770, n16256);
  not g30771 (n_14771, n16258);
  and g30772 (n16259, n_14770, n_14771);
  and g30773 (n16260, n5344, n7433);
  and g30774 (n16261, n6453, n10905);
  and g30775 (n16262, n5413, n7699);
  not g30776 (n_14772, n16261);
  not g30777 (n_14773, n16262);
  and g30778 (n16263, n_14772, n_14773);
  not g30779 (n_14774, n16260);
  not g30780 (n_14775, n16263);
  and g30781 (n16264, n_14774, n_14775);
  not g30782 (n_14776, n16264);
  and g30783 (n16265, \a[54] , n_14776);
  and g30784 (n16266, \a[40] , n16265);
  and g30785 (n16267, \a[42] , \a[52] );
  not g30786 (n_14777, n8239);
  not g30787 (n_14778, n16267);
  and g30788 (n16268, n_14777, n_14778);
  and g30789 (n16269, n_14774, n_14776);
  not g30790 (n_14779, n16268);
  and g30791 (n16270, n_14779, n16269);
  not g30792 (n_14780, n16266);
  not g30793 (n_14781, n16270);
  and g30794 (n16271, n_14780, n_14781);
  not g30795 (n_14782, n16259);
  not g30796 (n_14783, n16271);
  and g30797 (n16272, n_14782, n_14783);
  not g30798 (n_14784, n16272);
  and g30799 (n16273, n_14782, n_14784);
  and g30800 (n16274, n_14783, n_14784);
  not g30801 (n_14785, n16273);
  not g30802 (n_14786, n16274);
  and g30803 (n16275, n_14785, n_14786);
  and g30804 (n16276, n8503, n14569);
  and g30805 (n16277, n5560, n6256);
  not g30806 (n_14787, n16276);
  not g30807 (n_14788, n16277);
  and g30808 (n16278, n_14787, n_14788);
  and g30809 (n16279, n8578, n14569);
  not g30810 (n_14789, n16278);
  not g30811 (n_14790, n16279);
  and g30812 (n16280, n_14789, n_14790);
  not g30813 (n_14791, n16280);
  and g30814 (n16281, n8503, n_14791);
  and g30815 (n16282, n_14790, n_14791);
  not g30816 (n_14792, n8578);
  not g30817 (n_14793, n14569);
  and g30818 (n16283, n_14792, n_14793);
  not g30819 (n_14794, n16283);
  and g30820 (n16284, n16282, n_14794);
  not g30821 (n_14795, n16281);
  not g30822 (n_14796, n16284);
  and g30823 (n16285, n_14795, n_14796);
  not g30824 (n_14797, n16275);
  not g30825 (n_14798, n16285);
  and g30826 (n16286, n_14797, n_14798);
  not g30827 (n_14799, n16286);
  and g30828 (n16287, n_14797, n_14799);
  and g30829 (n16288, n_14798, n_14799);
  not g30830 (n_14800, n16287);
  not g30831 (n_14801, n16288);
  and g30832 (n16289, n_14800, n_14801);
  and g30833 (n16290, n_14604, n_14608);
  and g30834 (n16291, n16289, n16290);
  not g30835 (n_14802, n16289);
  not g30836 (n_14803, n16290);
  and g30837 (n16292, n_14802, n_14803);
  not g30838 (n_14804, n16291);
  not g30839 (n_14805, n16292);
  and g30840 (n16293, n_14804, n_14805);
  and g30841 (n16294, n2972, n8905);
  and g30842 (n16295, \a[59] , \a[62] );
  and g30843 (n16296, n6823, n16295);
  and g30844 (n16297, n3143, n9721);
  not g30845 (n_14806, n16296);
  not g30846 (n_14807, n16297);
  and g30847 (n16298, n_14806, n_14807);
  not g30848 (n_14808, n16294);
  not g30849 (n_14809, n16298);
  and g30850 (n16299, n_14808, n_14809);
  not g30851 (n_14810, n16299);
  and g30852 (n16300, \a[62] , n_14810);
  and g30853 (n16301, \a[32] , n16300);
  and g30854 (n16302, n_14808, n_14810);
  and g30855 (n16303, \a[33] , \a[61] );
  and g30856 (n16304, \a[35] , \a[59] );
  not g30857 (n_14811, n16303);
  not g30858 (n_14812, n16304);
  and g30859 (n16305, n_14811, n_14812);
  not g30860 (n_14813, n16305);
  and g30861 (n16306, n16302, n_14813);
  not g30862 (n_14814, n16301);
  not g30863 (n_14815, n16306);
  and g30864 (n16307, n_14814, n_14815);
  not g30865 (n_14816, n16307);
  and g30866 (n16308, n16185, n_14816);
  not g30867 (n_14817, n16185);
  and g30868 (n16309, n_14817, n16307);
  not g30869 (n_14818, n16308);
  not g30870 (n_14819, n16309);
  and g30871 (n16310, n_14818, n_14819);
  and g30872 (n16311, n5430, n11718);
  and g30873 (n16312, n11615, n13212);
  not g30874 (n_14820, n16311);
  not g30875 (n_14821, n16312);
  and g30876 (n16313, n_14820, n_14821);
  and g30877 (n16314, \a[34] , \a[60] );
  and g30878 (n16315, \a[39] , \a[55] );
  and g30879 (n16316, n16314, n16315);
  not g30880 (n_14822, n16313);
  not g30881 (n_14823, n16316);
  and g30882 (n16317, n_14822, n_14823);
  not g30883 (n_14824, n16317);
  and g30884 (n16318, \a[57] , n_14824);
  and g30885 (n16319, \a[37] , n16318);
  and g30886 (n16320, n_14823, n_14824);
  not g30887 (n_14825, n16314);
  not g30888 (n_14826, n16315);
  and g30889 (n16321, n_14825, n_14826);
  not g30890 (n_14827, n16321);
  and g30891 (n16322, n16320, n_14827);
  not g30892 (n_14828, n16319);
  not g30893 (n_14829, n16322);
  and g30894 (n16323, n_14828, n_14829);
  not g30895 (n_14830, n16310);
  not g30896 (n_14831, n16323);
  and g30897 (n16324, n_14830, n_14831);
  and g30898 (n16325, n16310, n16323);
  not g30899 (n_14832, n16324);
  not g30900 (n_14833, n16325);
  and g30901 (n16326, n_14832, n_14833);
  and g30902 (n16327, n16293, n16326);
  not g30903 (n_14834, n16293);
  not g30904 (n_14835, n16326);
  and g30905 (n16328, n_14834, n_14835);
  and g30906 (n16329, n_14611, n_14639);
  not g30907 (n_14836, n16198);
  and g30908 (n16330, n13038, n_14836);
  not g30909 (n_14837, n13038);
  and g30910 (n16331, n_14837, n16198);
  not g30911 (n_14838, n16330);
  not g30912 (n_14839, n16331);
  and g30913 (n16332, n_14838, n_14839);
  not g30914 (n_14840, n16332);
  and g30915 (n16333, n16173, n_14840);
  not g30916 (n_14841, n16173);
  and g30917 (n16334, n_14841, n16332);
  not g30918 (n_14842, n16333);
  not g30919 (n_14843, n16334);
  and g30920 (n16335, n_14842, n_14843);
  and g30921 (n16336, n_14704, n_14716);
  not g30922 (n_14844, n16335);
  and g30923 (n16337, n_14844, n16336);
  not g30924 (n_14845, n16336);
  and g30925 (n16338, n16335, n_14845);
  not g30926 (n_14846, n16337);
  not g30927 (n_14847, n16338);
  and g30928 (n16339, n_14846, n_14847);
  and g30929 (n16340, n16127, n16142);
  not g30930 (n_14848, n16127);
  not g30931 (n_14849, n16142);
  and g30932 (n16341, n_14848, n_14849);
  not g30933 (n_14850, n16340);
  not g30934 (n_14851, n16341);
  and g30935 (n16342, n_14850, n_14851);
  not g30936 (n_14852, n16342);
  and g30937 (n16343, n16158, n_14852);
  not g30938 (n_14853, n16158);
  and g30939 (n16344, n_14853, n16342);
  not g30940 (n_14854, n16343);
  not g30941 (n_14855, n16344);
  and g30942 (n16345, n_14854, n_14855);
  and g30943 (n16346, n16339, n16345);
  not g30944 (n_14856, n16339);
  not g30945 (n_14857, n16345);
  and g30946 (n16347, n_14856, n_14857);
  not g30947 (n_14858, n16346);
  not g30948 (n_14859, n16347);
  and g30949 (n16348, n_14858, n_14859);
  not g30950 (n_14860, n16329);
  and g30951 (n16349, n_14860, n16348);
  not g30952 (n_14861, n16348);
  and g30953 (n16350, n16329, n_14861);
  not g30954 (n_14862, n16349);
  not g30955 (n_14863, n16350);
  and g30956 (n16351, n_14862, n_14863);
  not g30957 (n_14864, n16328);
  and g30958 (n16352, n_14864, n16351);
  not g30959 (n_14865, n16327);
  and g30960 (n16353, n_14865, n16352);
  not g30961 (n_14866, n16353);
  and g30962 (n16354, n16351, n_14866);
  and g30963 (n16355, n_14864, n_14866);
  and g30964 (n16356, n_14865, n16355);
  not g30965 (n_14867, n16354);
  not g30966 (n_14868, n16356);
  and g30967 (n16357, n_14867, n_14868);
  not g30968 (n_14869, n16248);
  and g30969 (n16358, n_14869, n16357);
  not g30970 (n_14870, n16357);
  and g30971 (n16359, n16248, n_14870);
  not g30972 (n_14871, n16358);
  not g30973 (n_14872, n16359);
  and g30974 (n16360, n_14871, n_14872);
  and g30975 (n16361, n_14644, n_14737);
  not g30976 (n_14873, n16360);
  and g30977 (n16362, n_14873, n16361);
  not g30978 (n_14874, n16361);
  and g30979 (n16363, n16360, n_14874);
  not g30980 (n_14875, n16362);
  not g30981 (n_14876, n16363);
  and g30982 (n16364, n_14875, n_14876);
  and g30983 (n16365, n_14743, n_14742);
  not g30984 (n_14877, n16365);
  and g30985 (n16366, n_14741, n_14877);
  not g30986 (n_14878, n16364);
  and g30987 (n16367, n_14878, n16366);
  not g30988 (n_14879, n16366);
  and g30989 (n16368, n16364, n_14879);
  not g30990 (n_14880, n16367);
  not g30991 (n_14881, n16368);
  and g30992 (\asquared[95] , n_14880, n_14881);
  and g30993 (n16370, n_14862, n_14866);
  and g30994 (n16371, n_14805, n_14865);
  and g30995 (n16372, n3828, n9509);
  not g30996 (n_14882, n16372);
  and g30997 (n16373, \a[59] , n_14882);
  and g30998 (n16374, \a[36] , n16373);
  and g30999 (n16375, \a[60] , n_14882);
  and g31000 (n16376, \a[35] , n16375);
  not g31001 (n_14883, n16374);
  not g31002 (n_14884, n16376);
  and g31003 (n16377, n_14883, n_14884);
  not g31004 (n_14885, n16282);
  not g31005 (n_14886, n16377);
  and g31006 (n16378, n_14885, n_14886);
  not g31007 (n_14887, n16378);
  and g31008 (n16379, n_14885, n_14887);
  and g31009 (n16380, n_14886, n_14887);
  not g31010 (n_14888, n16379);
  not g31011 (n_14889, n16380);
  and g31012 (n16381, n_14888, n_14889);
  and g31013 (n16382, n_14838, n_14843);
  and g31014 (n16383, n16381, n16382);
  not g31015 (n_14890, n16381);
  not g31016 (n_14891, n16382);
  and g31017 (n16384, n_14890, n_14891);
  not g31018 (n_14892, n16383);
  not g31019 (n_14893, n16384);
  and g31020 (n16385, n_14892, n_14893);
  and g31021 (n16386, n_14851, n_14855);
  not g31022 (n_14894, n16385);
  and g31023 (n16387, n_14894, n16386);
  not g31024 (n_14895, n16386);
  and g31025 (n16388, n16385, n_14895);
  not g31026 (n_14896, n16387);
  not g31027 (n_14897, n16388);
  and g31028 (n16389, n_14896, n_14897);
  and g31029 (n16390, n_14847, n_14858);
  not g31030 (n_14898, n16390);
  and g31031 (n16391, n16389, n_14898);
  not g31032 (n_14899, n16389);
  and g31033 (n16392, n_14899, n16390);
  not g31034 (n_14900, n16391);
  not g31035 (n_14901, n16392);
  and g31036 (n16393, n_14900, n_14901);
  not g31037 (n_14902, n16371);
  and g31038 (n16394, n_14902, n16393);
  not g31039 (n_14903, n16393);
  and g31040 (n16395, n16371, n_14903);
  not g31041 (n_14904, n16394);
  not g31042 (n_14905, n16395);
  and g31043 (n16396, n_14904, n_14905);
  not g31044 (n_14906, n16396);
  and g31045 (n16397, n16370, n_14906);
  not g31046 (n_14907, n16370);
  and g31047 (n16398, n_14907, n16396);
  not g31048 (n_14908, n16397);
  not g31049 (n_14909, n16398);
  and g31050 (n16399, n_14908, n_14909);
  and g31051 (n16400, \a[48] , \a[62] );
  and g31052 (n16401, \a[33] , n16400);
  not g31053 (n_14910, n16401);
  and g31054 (n16402, n6252, n_14910);
  not g31055 (n_14911, n16402);
  and g31056 (n16403, n_14910, n_14911);
  and g31057 (n16404, \a[33] , \a[62] );
  not g31058 (n_14912, \a[48] );
  not g31059 (n_14913, n16404);
  and g31060 (n16405, n_14912, n_14913);
  not g31061 (n_14914, n16405);
  and g31062 (n16406, n16403, n_14914);
  and g31063 (n16407, n6252, n_14911);
  not g31064 (n_14915, n16406);
  not g31065 (n_14916, n16407);
  and g31066 (n16408, n_14915, n_14916);
  and g31067 (n16409, n5560, n6325);
  and g31068 (n16410, \a[46] , \a[49] );
  not g31069 (n_14917, n8506);
  not g31070 (n_14918, n16410);
  and g31071 (n16411, n_14917, n_14918);
  not g31072 (n_14919, n16409);
  not g31073 (n_14920, n16411);
  not g31077 (n_14921, n16414);
  and g31078 (n16415, \a[56] , n_14921);
  and g31079 (n16416, \a[39] , n16415);
  and g31080 (n16417, n_14919, n_14921);
  and g31081 (n16418, n_14920, n16417);
  not g31082 (n_14922, n16416);
  not g31083 (n_14923, n16418);
  and g31084 (n16419, n_14922, n_14923);
  not g31085 (n_14924, n16408);
  not g31086 (n_14925, n16419);
  and g31087 (n16420, n_14924, n_14925);
  not g31088 (n_14926, n16420);
  and g31089 (n16421, n_14924, n_14926);
  and g31090 (n16422, n_14925, n_14926);
  not g31091 (n_14927, n16421);
  not g31092 (n_14928, n16422);
  and g31093 (n16423, n_14927, n_14928);
  and g31094 (n16424, n5296, n6968);
  and g31095 (n16425, n4639, n7232);
  and g31096 (n16426, n5018, n7433);
  not g31097 (n_14929, n16425);
  not g31098 (n_14930, n16426);
  and g31099 (n16427, n_14929, n_14930);
  not g31100 (n_14931, n16424);
  not g31101 (n_14932, n16427);
  and g31102 (n16428, n_14931, n_14932);
  not g31103 (n_14933, n16428);
  and g31104 (n16429, \a[53] , n_14933);
  and g31105 (n16430, \a[42] , n16429);
  and g31106 (n16431, \a[43] , \a[52] );
  not g31107 (n_14934, n8486);
  not g31108 (n_14935, n16431);
  and g31109 (n16432, n_14934, n_14935);
  and g31110 (n16433, n_14931, n_14933);
  not g31111 (n_14936, n16432);
  and g31112 (n16434, n_14936, n16433);
  not g31113 (n_14937, n16430);
  not g31114 (n_14938, n16434);
  and g31115 (n16435, n_14937, n_14938);
  not g31116 (n_14939, n16423);
  not g31117 (n_14940, n16435);
  and g31118 (n16436, n_14939, n_14940);
  not g31119 (n_14941, n16436);
  and g31120 (n16437, n_14939, n_14941);
  and g31121 (n16438, n_14940, n_14941);
  not g31122 (n_14942, n16437);
  not g31123 (n_14943, n16438);
  and g31124 (n16439, n_14942, n_14943);
  and g31125 (n16440, n_14748, n_14752);
  and g31126 (n16441, n16439, n16440);
  not g31127 (n_14944, n16439);
  not g31128 (n_14945, n16440);
  and g31129 (n16442, n_14944, n_14945);
  not g31130 (n_14946, n16441);
  not g31131 (n_14947, n16442);
  and g31132 (n16443, n_14946, n_14947);
  and g31133 (n16444, \a[32] , \a[63] );
  and g31134 (n16445, \a[34] , \a[61] );
  not g31135 (n_14948, n16444);
  not g31136 (n_14949, n16445);
  and g31137 (n16446, n_14948, n_14949);
  and g31138 (n16447, n4090, n9909);
  not g31139 (n_14950, n16447);
  not g31142 (n_14951, n16446);
  not g31144 (n_14952, n16450);
  and g31145 (n16451, n_14950, n_14952);
  and g31146 (n16452, n_14951, n16451);
  and g31147 (n16453, \a[54] , n_14952);
  and g31148 (n16454, \a[41] , n16453);
  not g31149 (n_14953, n16452);
  not g31150 (n_14954, n16454);
  and g31151 (n16455, n_14953, n_14954);
  and g31152 (n16456, n3803, n11718);
  and g31153 (n16457, \a[55] , \a[58] );
  and g31154 (n16458, n5695, n16457);
  and g31155 (n16459, n4565, n8436);
  not g31156 (n_14955, n16458);
  not g31157 (n_14956, n16459);
  and g31158 (n16460, n_14955, n_14956);
  not g31159 (n_14957, n16456);
  not g31160 (n_14958, n16460);
  and g31161 (n16461, n_14957, n_14958);
  not g31162 (n_14959, n16461);
  and g31163 (n16462, \a[37] , n_14959);
  and g31164 (n16463, \a[58] , n16462);
  and g31165 (n16464, n_14957, n_14959);
  and g31166 (n16465, \a[38] , \a[57] );
  and g31167 (n16466, \a[40] , \a[55] );
  not g31168 (n_14960, n16465);
  not g31169 (n_14961, n16466);
  and g31170 (n16467, n_14960, n_14961);
  not g31171 (n_14962, n16467);
  and g31172 (n16468, n16464, n_14962);
  not g31173 (n_14963, n16463);
  not g31174 (n_14964, n16468);
  and g31175 (n16469, n_14963, n_14964);
  not g31176 (n_14965, n16255);
  not g31177 (n_14966, n16469);
  and g31178 (n16470, n_14965, n_14966);
  not g31179 (n_14967, n16470);
  and g31180 (n16471, n_14965, n_14967);
  and g31181 (n16472, n_14966, n_14967);
  not g31182 (n_14968, n16471);
  not g31183 (n_14969, n16472);
  and g31184 (n16473, n_14968, n_14969);
  not g31185 (n_14970, n16455);
  not g31186 (n_14971, n16473);
  and g31187 (n16474, n_14970, n_14971);
  not g31188 (n_14972, n16474);
  and g31189 (n16475, n_14970, n_14972);
  and g31190 (n16476, n_14971, n_14972);
  not g31191 (n_14973, n16475);
  not g31192 (n_14974, n16476);
  and g31193 (n16477, n_14973, n_14974);
  not g31194 (n_14975, n16477);
  and g31195 (n16478, n16443, n_14975);
  not g31196 (n_14976, n16478);
  and g31197 (n16479, n16443, n_14976);
  and g31198 (n16480, n_14975, n_14976);
  not g31199 (n_14977, n16479);
  not g31200 (n_14978, n16480);
  and g31201 (n16481, n_14977, n_14978);
  and g31202 (n16482, n_14755, n_14759);
  and g31203 (n16483, n16302, n16320);
  not g31204 (n_14979, n16302);
  not g31205 (n_14980, n16320);
  and g31206 (n16484, n_14979, n_14980);
  not g31207 (n_14981, n16483);
  not g31208 (n_14982, n16484);
  and g31209 (n16485, n_14981, n_14982);
  not g31210 (n_14983, n16485);
  and g31211 (n16486, n16269, n_14983);
  not g31212 (n_14984, n16269);
  and g31213 (n16487, n_14984, n16485);
  not g31214 (n_14985, n16486);
  not g31215 (n_14986, n16487);
  and g31216 (n16488, n_14985, n_14986);
  and g31217 (n16489, n_14784, n_14799);
  and g31218 (n16490, n_14817, n_14816);
  not g31219 (n_14987, n16490);
  and g31220 (n16491, n_14832, n_14987);
  and g31221 (n16492, n16489, n16491);
  not g31222 (n_14988, n16489);
  not g31223 (n_14989, n16491);
  and g31224 (n16493, n_14988, n_14989);
  not g31225 (n_14990, n16492);
  not g31226 (n_14991, n16493);
  and g31227 (n16494, n_14990, n_14991);
  and g31228 (n16495, n16488, n16494);
  not g31229 (n_14992, n16488);
  not g31230 (n_14993, n16494);
  and g31231 (n16496, n_14992, n_14993);
  not g31232 (n_14994, n16495);
  not g31233 (n_14995, n16496);
  and g31234 (n16497, n_14994, n_14995);
  not g31235 (n_14996, n16482);
  and g31236 (n16498, n_14996, n16497);
  not g31237 (n_14997, n16497);
  and g31238 (n16499, n16482, n_14997);
  not g31239 (n_14998, n16498);
  not g31240 (n_14999, n16499);
  and g31241 (n16500, n_14998, n_14999);
  and g31242 (n16501, n16481, n16500);
  not g31243 (n_15000, n16481);
  not g31244 (n_15001, n16500);
  and g31245 (n16502, n_15000, n_15001);
  not g31246 (n_15002, n16501);
  not g31247 (n_15003, n16502);
  and g31248 (n16503, n_15002, n_15003);
  not g31249 (n_15004, n16503);
  and g31250 (n16504, n16399, n_15004);
  not g31251 (n_15005, n16504);
  and g31252 (n16505, n16399, n_15005);
  and g31253 (n16506, n_15004, n_15005);
  not g31254 (n_15006, n16505);
  not g31255 (n_15007, n16506);
  and g31256 (n16507, n_15006, n_15007);
  and g31257 (n16508, n_14764, n_14872);
  not g31258 (n_15008, n16507);
  not g31259 (n_15009, n16508);
  and g31260 (n16509, n_15008, n_15009);
  and g31261 (n16510, n16507, n16508);
  not g31262 (n_15010, n16509);
  not g31263 (n_15011, n16510);
  and g31264 (n16511, n_15010, n_15011);
  and g31265 (n16512, n_14875, n_14879);
  not g31266 (n_15012, n16512);
  and g31267 (n16513, n_14876, n_15012);
  not g31268 (n_15013, n16511);
  and g31269 (n16514, n_15013, n16513);
  not g31270 (n_15014, n16513);
  and g31271 (n16515, n16511, n_15014);
  not g31272 (n_15015, n16514);
  not g31273 (n_15016, n16515);
  and g31274 (\asquared[96] , n_15015, n_15016);
  and g31275 (n16517, n_15011, n_15014);
  not g31276 (n_15017, n16517);
  and g31277 (n16518, n_15010, n_15017);
  and g31278 (n16519, n_14909, n_15005);
  and g31279 (n16520, n_14947, n_14976);
  and g31280 (n16521, n5695, n13870);
  and g31281 (n16522, n3687, n9509);
  and g31282 (n16523, \a[40] , \a[60] );
  and g31283 (n16524, n15987, n16523);
  not g31284 (n_15018, n16522);
  not g31285 (n_15019, n16524);
  and g31286 (n16525, n_15018, n_15019);
  not g31287 (n_15020, n16521);
  not g31288 (n_15021, n16525);
  and g31289 (n16526, n_15020, n_15021);
  not g31290 (n_15022, n16526);
  and g31291 (n16527, n_15020, n_15022);
  and g31292 (n16528, \a[37] , \a[59] );
  and g31293 (n16529, \a[40] , \a[56] );
  not g31294 (n_15023, n16528);
  not g31295 (n_15024, n16529);
  and g31296 (n16530, n_15023, n_15024);
  not g31297 (n_15025, n16530);
  and g31298 (n16531, n16527, n_15025);
  and g31299 (n16532, \a[60] , n_15022);
  and g31300 (n16533, \a[36] , n16532);
  not g31301 (n_15026, n16531);
  not g31302 (n_15027, n16533);
  and g31303 (n16534, n_15026, n_15027);
  and g31304 (n16535, \a[38] , \a[58] );
  and g31305 (n16536, \a[39] , \a[57] );
  not g31306 (n_15028, n16535);
  not g31307 (n_15029, n16536);
  and g31308 (n16537, n_15028, n_15029);
  and g31309 (n16538, n5083, n8436);
  not g31310 (n_15030, n16538);
  and g31311 (n16539, n8700, n_15030);
  not g31312 (n_15031, n16537);
  and g31313 (n16540, n_15031, n16539);
  not g31314 (n_15032, n16540);
  and g31315 (n16541, n8700, n_15032);
  and g31316 (n16542, n_15030, n_15032);
  and g31317 (n16543, n_15031, n16542);
  not g31318 (n_15033, n16541);
  not g31319 (n_15034, n16543);
  and g31320 (n16544, n_15033, n_15034);
  not g31321 (n_15035, n16534);
  not g31322 (n_15036, n16544);
  and g31323 (n16545, n_15035, n_15036);
  not g31324 (n_15037, n16545);
  and g31325 (n16546, n_15035, n_15037);
  and g31326 (n16547, n_15036, n_15037);
  not g31327 (n_15038, n16546);
  not g31328 (n_15039, n16547);
  and g31329 (n16548, n_15038, n_15039);
  and g31330 (n16549, \a[45] , \a[51] );
  and g31331 (n16550, n5666, n6325);
  and g31332 (n16551, n6254, n16549);
  and g31333 (n16552, n5560, n6564);
  not g31334 (n_15040, n16551);
  not g31335 (n_15041, n16552);
  and g31336 (n16553, n_15040, n_15041);
  not g31337 (n_15042, n16550);
  not g31338 (n_15043, n16553);
  and g31339 (n16554, n_15042, n_15043);
  not g31340 (n_15044, n16554);
  and g31341 (n16555, n16549, n_15044);
  and g31342 (n16556, n_15042, n_15044);
  and g31343 (n16557, \a[46] , \a[50] );
  not g31344 (n_15045, n6254);
  not g31345 (n_15046, n16557);
  and g31346 (n16558, n_15045, n_15046);
  not g31347 (n_15047, n16558);
  and g31348 (n16559, n16556, n_15047);
  not g31349 (n_15048, n16555);
  not g31350 (n_15049, n16559);
  and g31351 (n16560, n_15048, n_15049);
  not g31352 (n_15050, n16548);
  not g31353 (n_15051, n16560);
  and g31354 (n16561, n_15050, n_15051);
  not g31355 (n_15052, n16561);
  and g31356 (n16562, n_15050, n_15052);
  and g31357 (n16563, n_15051, n_15052);
  not g31358 (n_15053, n16562);
  not g31359 (n_15054, n16563);
  and g31360 (n16564, n_15053, n_15054);
  and g31361 (n16565, n_14991, n_14994);
  not g31362 (n_15055, n16564);
  not g31363 (n_15056, n16565);
  and g31364 (n16566, n_15055, n_15056);
  not g31365 (n_15057, n16566);
  and g31366 (n16567, n_15055, n_15057);
  and g31367 (n16568, n_15056, n_15057);
  not g31368 (n_15058, n16567);
  not g31369 (n_15059, n16568);
  and g31370 (n16569, n_15058, n_15059);
  not g31371 (n_15060, n16520);
  not g31372 (n_15061, n16569);
  and g31373 (n16570, n_15060, n_15061);
  not g31374 (n_15062, n16570);
  and g31375 (n16571, n_15060, n_15062);
  and g31376 (n16572, n_15061, n_15062);
  not g31377 (n_15063, n16571);
  not g31378 (n_15064, n16572);
  and g31379 (n16573, n_15063, n_15064);
  and g31380 (n16574, n_15000, n16500);
  not g31381 (n_15065, n16574);
  and g31382 (n16575, n_14998, n_15065);
  not g31383 (n_15066, n16573);
  not g31384 (n_15067, n16575);
  and g31385 (n16576, n_15066, n_15067);
  not g31386 (n_15068, n16576);
  and g31387 (n16577, n_15066, n_15068);
  and g31388 (n16578, n_15067, n_15068);
  not g31389 (n_15069, n16577);
  not g31390 (n_15070, n16578);
  and g31391 (n16579, n_15069, n_15070);
  and g31392 (n16580, n_14900, n_14904);
  and g31393 (n16581, n16403, n16417);
  not g31394 (n_15071, n16403);
  not g31395 (n_15072, n16417);
  and g31396 (n16582, n_15071, n_15072);
  not g31397 (n_15073, n16581);
  not g31398 (n_15074, n16582);
  and g31399 (n16583, n_15073, n_15074);
  not g31400 (n_15075, n16583);
  and g31401 (n16584, n16433, n_15075);
  not g31402 (n_15076, n16433);
  and g31403 (n16585, n_15076, n16583);
  not g31404 (n_15077, n16584);
  not g31405 (n_15078, n16585);
  and g31406 (n16586, n_15077, n_15078);
  and g31407 (n16587, n_14967, n_14972);
  and g31408 (n16588, n_14926, n_14941);
  and g31409 (n16589, n16587, n16588);
  not g31410 (n_15079, n16587);
  not g31411 (n_15080, n16588);
  and g31412 (n16590, n_15079, n_15080);
  not g31413 (n_15081, n16589);
  not g31414 (n_15082, n16590);
  and g31415 (n16591, n_15081, n_15082);
  and g31416 (n16592, n16586, n16591);
  not g31417 (n_15083, n16586);
  not g31418 (n_15084, n16591);
  and g31419 (n16593, n_15083, n_15084);
  not g31420 (n_15085, n16592);
  not g31421 (n_15086, n16593);
  and g31422 (n16594, n_15085, n_15086);
  not g31423 (n_15087, n16580);
  and g31424 (n16595, n_15087, n16594);
  not g31425 (n_15088, n16594);
  and g31426 (n16596, n16580, n_15088);
  not g31427 (n_15089, n16595);
  not g31428 (n_15090, n16596);
  and g31429 (n16597, n_15089, n_15090);
  and g31430 (n16598, n3319, n9721);
  and g31431 (n16599, n2972, n9909);
  and g31432 (n16600, n4150, n9792);
  not g31433 (n_15091, n16599);
  not g31434 (n_15092, n16600);
  and g31435 (n16601, n_15091, n_15092);
  not g31436 (n_15093, n16598);
  not g31437 (n_15094, n16601);
  and g31438 (n16602, n_15093, n_15094);
  not g31439 (n_15095, n16602);
  and g31440 (n16603, n_15093, n_15095);
  and g31441 (n16604, \a[34] , \a[62] );
  and g31442 (n16605, \a[35] , \a[61] );
  not g31443 (n_15096, n16604);
  not g31444 (n_15097, n16605);
  and g31445 (n16606, n_15096, n_15097);
  not g31446 (n_15098, n16606);
  and g31447 (n16607, n16603, n_15098);
  and g31448 (n16608, \a[63] , n_15095);
  and g31449 (n16609, \a[33] , n16608);
  not g31450 (n_15099, n16607);
  not g31451 (n_15100, n16609);
  and g31452 (n16610, n_15099, n_15100);
  and g31453 (n16611, n5018, n7699);
  and g31454 (n16612, \a[43] , \a[53] );
  and g31455 (n16613, n8594, n16612);
  and g31456 (n16614, n5344, n7701);
  not g31457 (n_15101, n16613);
  not g31458 (n_15102, n16614);
  and g31459 (n16615, n_15101, n_15102);
  not g31460 (n_15103, n16611);
  not g31461 (n_15104, n16615);
  and g31462 (n16616, n_15103, n_15104);
  not g31463 (n_15105, n16616);
  and g31464 (n16617, n8594, n_15105);
  and g31465 (n16618, \a[42] , \a[54] );
  not g31466 (n_15106, n16612);
  not g31467 (n_15107, n16618);
  and g31468 (n16619, n_15106, n_15107);
  and g31469 (n16620, n_15103, n_15105);
  not g31470 (n_15108, n16619);
  and g31471 (n16621, n_15108, n16620);
  not g31472 (n_15109, n16617);
  not g31473 (n_15110, n16621);
  and g31474 (n16622, n_15109, n_15110);
  not g31475 (n_15111, n16610);
  not g31476 (n_15112, n16622);
  and g31477 (n16623, n_15111, n_15112);
  not g31478 (n_15113, n16623);
  and g31479 (n16624, n_15111, n_15113);
  and g31480 (n16625, n_15112, n_15113);
  not g31481 (n_15114, n16624);
  not g31482 (n_15115, n16625);
  and g31483 (n16626, n_15114, n_15115);
  and g31484 (n16627, n_14982, n_14986);
  and g31485 (n16628, n16626, n16627);
  not g31486 (n_15116, n16626);
  not g31487 (n_15117, n16627);
  and g31488 (n16629, n_15116, n_15117);
  not g31489 (n_15118, n16628);
  not g31490 (n_15119, n16629);
  and g31491 (n16630, n_15118, n_15119);
  and g31492 (n16631, n16451, n16464);
  not g31493 (n_15120, n16451);
  not g31494 (n_15121, n16464);
  and g31495 (n16632, n_15120, n_15121);
  not g31496 (n_15122, n16631);
  not g31497 (n_15123, n16632);
  and g31498 (n16633, n_15122, n_15123);
  and g31499 (n16634, n_14882, n_14887);
  not g31500 (n_15124, n16633);
  and g31501 (n16635, n_15124, n16634);
  not g31502 (n_15125, n16634);
  and g31503 (n16636, n16633, n_15125);
  not g31504 (n_15126, n16635);
  not g31505 (n_15127, n16636);
  and g31506 (n16637, n_15126, n_15127);
  and g31507 (n16638, n_14893, n_14897);
  not g31508 (n_15128, n16637);
  and g31509 (n16639, n_15128, n16638);
  not g31510 (n_15129, n16638);
  and g31511 (n16640, n16637, n_15129);
  not g31512 (n_15130, n16639);
  not g31513 (n_15131, n16640);
  and g31514 (n16641, n_15130, n_15131);
  and g31515 (n16642, n16630, n16641);
  not g31516 (n_15132, n16630);
  not g31517 (n_15133, n16641);
  and g31518 (n16643, n_15132, n_15133);
  not g31519 (n_15134, n16642);
  not g31520 (n_15135, n16643);
  and g31521 (n16644, n_15134, n_15135);
  and g31522 (n16645, n16597, n16644);
  not g31523 (n_15136, n16597);
  not g31524 (n_15137, n16644);
  and g31525 (n16646, n_15136, n_15137);
  not g31526 (n_15138, n16645);
  not g31527 (n_15139, n16646);
  and g31528 (n16647, n_15138, n_15139);
  not g31529 (n_15140, n16579);
  and g31530 (n16648, n_15140, n16647);
  not g31531 (n_15141, n16647);
  and g31532 (n16649, n_15070, n_15141);
  and g31533 (n16650, n_15069, n16649);
  not g31534 (n_15142, n16648);
  not g31535 (n_15143, n16650);
  and g31536 (n16651, n_15142, n_15143);
  not g31537 (n_15144, n16651);
  and g31538 (n16652, n16519, n_15144);
  not g31539 (n_15145, n16519);
  and g31540 (n16653, n_15145, n16651);
  not g31541 (n_15146, n16652);
  not g31542 (n_15147, n16653);
  and g31543 (n16654, n_15146, n_15147);
  not g31544 (n_15148, n16654);
  and g31545 (n16655, n16518, n_15148);
  not g31546 (n_15149, n16518);
  and g31547 (n16656, n_15149, n_15146);
  and g31548 (n16657, n_15147, n16656);
  not g31549 (n_15150, n16655);
  not g31550 (n_15151, n16657);
  and g31551 (\asquared[97] , n_15150, n_15151);
  not g31552 (n_15152, n16656);
  and g31553 (n16659, n_15147, n_15152);
  and g31554 (n16660, n_15068, n_15142);
  and g31555 (n16661, n_15057, n_15062);
  and g31556 (n16662, \a[36] , \a[61] );
  not g31557 (n_15153, n16556);
  and g31558 (n16663, n_15153, n16662);
  not g31559 (n_15154, n16662);
  and g31560 (n16664, n16556, n_15154);
  not g31561 (n_15155, n16663);
  not g31562 (n_15156, n16664);
  and g31563 (n16665, n_15155, n_15156);
  not g31564 (n_15157, n16665);
  and g31565 (n16666, n16542, n_15157);
  not g31566 (n_15158, n16542);
  and g31567 (n16667, n_15158, n16665);
  not g31568 (n_15159, n16666);
  not g31569 (n_15160, n16667);
  and g31570 (n16668, n_15159, n_15160);
  and g31571 (n16669, n_15037, n_15052);
  and g31572 (n16670, n_15123, n_15127);
  and g31573 (n16671, n16669, n16670);
  not g31574 (n_15161, n16669);
  not g31575 (n_15162, n16670);
  and g31576 (n16672, n_15161, n_15162);
  not g31577 (n_15163, n16671);
  not g31578 (n_15164, n16672);
  and g31579 (n16673, n_15163, n_15164);
  and g31580 (n16674, n16668, n16673);
  not g31581 (n_15165, n16668);
  not g31582 (n_15166, n16673);
  and g31583 (n16675, n_15165, n_15166);
  not g31584 (n_15167, n16674);
  not g31585 (n_15168, n16675);
  and g31586 (n16676, n_15167, n_15168);
  and g31587 (n16677, \a[49] , \a[62] );
  and g31588 (n16678, \a[35] , n16677);
  not g31589 (n_15169, n16678);
  and g31590 (n16679, n6256, n_15169);
  not g31591 (n_15170, n16679);
  and g31592 (n16680, n_15169, n_15170);
  and g31593 (n16681, \a[35] , \a[62] );
  not g31594 (n_15171, \a[49] );
  not g31595 (n_15172, n16681);
  and g31596 (n16682, n_15171, n_15172);
  not g31597 (n_15173, n16682);
  and g31598 (n16683, n16680, n_15173);
  and g31599 (n16684, n6256, n_15170);
  not g31600 (n_15174, n16683);
  not g31601 (n_15175, n16684);
  and g31602 (n16685, n_15174, n_15175);
  and g31603 (n16686, \a[47] , \a[50] );
  not g31604 (n_15176, n8854);
  not g31605 (n_15177, n16686);
  and g31606 (n16687, n_15176, n_15177);
  and g31607 (n16688, n5666, n6564);
  not g31608 (n_15178, n16688);
  not g31611 (n_15179, n16687);
  not g31613 (n_15180, n16691);
  and g31614 (n16692, \a[57] , n_15180);
  and g31615 (n16693, \a[40] , n16692);
  and g31616 (n16694, n_15178, n_15180);
  and g31617 (n16695, n_15179, n16694);
  not g31618 (n_15181, n16693);
  not g31619 (n_15182, n16695);
  and g31620 (n16696, n_15181, n_15182);
  not g31621 (n_15183, n16685);
  not g31622 (n_15184, n16696);
  and g31623 (n16697, n_15183, n_15184);
  not g31624 (n_15185, n16697);
  and g31625 (n16698, n_15183, n_15185);
  and g31626 (n16699, n_15184, n_15185);
  not g31627 (n_15186, n16698);
  not g31628 (n_15187, n16699);
  and g31629 (n16700, n_15186, n_15187);
  and g31630 (n16701, n_15074, n_15078);
  and g31631 (n16702, n16700, n16701);
  not g31632 (n_15188, n16700);
  not g31633 (n_15189, n16701);
  and g31634 (n16703, n_15188, n_15189);
  not g31635 (n_15190, n16702);
  not g31636 (n_15191, n16703);
  and g31637 (n16704, n_15190, n_15191);
  and g31638 (n16705, n16527, n16603);
  not g31639 (n_15192, n16527);
  not g31640 (n_15193, n16603);
  and g31641 (n16706, n_15192, n_15193);
  not g31642 (n_15194, n16705);
  not g31643 (n_15195, n16706);
  and g31644 (n16707, n_15194, n_15195);
  not g31645 (n_15196, n16707);
  and g31646 (n16708, n16620, n_15196);
  not g31647 (n_15197, n16620);
  and g31648 (n16709, n_15197, n16707);
  not g31649 (n_15198, n16708);
  not g31650 (n_15199, n16709);
  and g31651 (n16710, n_15198, n_15199);
  and g31652 (n16711, n_15113, n_15119);
  not g31653 (n_15200, n16710);
  and g31654 (n16712, n_15200, n16711);
  not g31655 (n_15201, n16711);
  and g31656 (n16713, n16710, n_15201);
  not g31657 (n_15202, n16712);
  not g31658 (n_15203, n16713);
  and g31659 (n16714, n_15202, n_15203);
  and g31660 (n16715, n16704, n16714);
  not g31661 (n_15204, n16704);
  not g31662 (n_15205, n16714);
  and g31663 (n16716, n_15204, n_15205);
  not g31664 (n_15206, n16715);
  not g31665 (n_15207, n16716);
  and g31666 (n16717, n_15206, n_15207);
  and g31667 (n16718, n16676, n16717);
  not g31668 (n_15208, n16676);
  not g31669 (n_15209, n16717);
  and g31670 (n16719, n_15208, n_15209);
  not g31671 (n_15210, n16718);
  not g31672 (n_15211, n16719);
  and g31673 (n16720, n_15210, n_15211);
  not g31674 (n_15212, n16720);
  and g31675 (n16721, n16661, n_15212);
  not g31676 (n_15213, n16661);
  and g31677 (n16722, n_15213, n16720);
  not g31678 (n_15214, n16721);
  not g31679 (n_15215, n16722);
  and g31680 (n16723, n_15214, n_15215);
  and g31681 (n16724, n_15131, n_15134);
  and g31682 (n16725, n5344, n9161);
  and g31683 (n16726, \a[34] , \a[63] );
  and g31684 (n16727, \a[41] , \a[56] );
  and g31685 (n16728, n16726, n16727);
  not g31686 (n_15216, n16725);
  not g31687 (n_15217, n16728);
  and g31688 (n16729, n_15216, n_15217);
  and g31689 (n16730, \a[42] , \a[55] );
  and g31690 (n16731, n16726, n16730);
  not g31691 (n_15218, n16729);
  not g31692 (n_15219, n16731);
  and g31693 (n16732, n_15218, n_15219);
  not g31694 (n_15220, n16732);
  and g31695 (n16733, n_15219, n_15220);
  not g31696 (n_15221, n16726);
  not g31697 (n_15222, n16730);
  and g31698 (n16734, n_15221, n_15222);
  not g31699 (n_15223, n16734);
  and g31700 (n16735, n16733, n_15223);
  and g31701 (n16736, n16727, n_15220);
  not g31702 (n_15224, n16735);
  not g31703 (n_15225, n16736);
  and g31704 (n16737, n_15224, n_15225);
  and g31705 (n16738, n5083, n8987);
  and g31706 (n16739, n5430, n10089);
  and g31707 (n16740, n4565, n9509);
  not g31708 (n_15226, n16739);
  not g31709 (n_15227, n16740);
  and g31710 (n16741, n_15226, n_15227);
  not g31711 (n_15228, n16738);
  not g31712 (n_15229, n16741);
  and g31713 (n16742, n_15228, n_15229);
  not g31714 (n_15230, n16742);
  and g31715 (n16743, \a[60] , n_15230);
  and g31716 (n16744, \a[37] , n16743);
  and g31717 (n16745, n_15228, n_15230);
  and g31718 (n16746, \a[38] , \a[59] );
  and g31719 (n16747, \a[39] , \a[58] );
  not g31720 (n_15231, n16746);
  not g31721 (n_15232, n16747);
  and g31722 (n16748, n_15231, n_15232);
  not g31723 (n_15233, n16748);
  and g31724 (n16749, n16745, n_15233);
  not g31725 (n_15234, n16744);
  not g31726 (n_15235, n16749);
  and g31727 (n16750, n_15234, n_15235);
  not g31728 (n_15236, n16737);
  not g31729 (n_15237, n16750);
  and g31730 (n16751, n_15236, n_15237);
  not g31731 (n_15238, n16751);
  and g31732 (n16752, n_15236, n_15238);
  and g31733 (n16753, n_15237, n_15238);
  not g31734 (n_15239, n16752);
  not g31735 (n_15240, n16753);
  and g31736 (n16754, n_15239, n_15240);
  and g31737 (n16755, n5713, n7433);
  and g31738 (n16756, n4811, n10905);
  and g31739 (n16757, n5296, n7699);
  not g31740 (n_15241, n16756);
  not g31741 (n_15242, n16757);
  and g31742 (n16758, n_15241, n_15242);
  not g31743 (n_15243, n16755);
  not g31744 (n_15244, n16758);
  and g31745 (n16759, n_15243, n_15244);
  not g31746 (n_15245, n16759);
  and g31747 (n16760, \a[54] , n_15245);
  and g31748 (n16761, \a[43] , n16760);
  and g31749 (n16762, \a[44] , \a[53] );
  not g31750 (n_15246, n9108);
  not g31751 (n_15247, n16762);
  and g31752 (n16763, n_15246, n_15247);
  and g31753 (n16764, n_15243, n_15245);
  not g31754 (n_15248, n16763);
  and g31755 (n16765, n_15248, n16764);
  not g31756 (n_15249, n16761);
  not g31757 (n_15250, n16765);
  and g31758 (n16766, n_15249, n_15250);
  not g31759 (n_15251, n16754);
  not g31760 (n_15252, n16766);
  and g31761 (n16767, n_15251, n_15252);
  not g31762 (n_15253, n16767);
  and g31763 (n16768, n_15251, n_15253);
  and g31764 (n16769, n_15252, n_15253);
  not g31765 (n_15254, n16768);
  not g31766 (n_15255, n16769);
  and g31767 (n16770, n_15254, n_15255);
  and g31768 (n16771, n_15082, n_15085);
  not g31769 (n_15256, n16770);
  not g31770 (n_15257, n16771);
  and g31771 (n16772, n_15256, n_15257);
  not g31772 (n_15258, n16772);
  and g31773 (n16773, n_15256, n_15258);
  and g31774 (n16774, n_15257, n_15258);
  not g31775 (n_15259, n16773);
  not g31776 (n_15260, n16774);
  and g31777 (n16775, n_15259, n_15260);
  not g31778 (n_15261, n16724);
  not g31779 (n_15262, n16775);
  and g31780 (n16776, n_15261, n_15262);
  not g31781 (n_15263, n16776);
  and g31782 (n16777, n_15261, n_15263);
  and g31783 (n16778, n_15262, n_15263);
  not g31784 (n_15264, n16777);
  not g31785 (n_15265, n16778);
  and g31786 (n16779, n_15264, n_15265);
  and g31787 (n16780, n_15089, n_15138);
  and g31788 (n16781, n16779, n16780);
  not g31789 (n_15266, n16779);
  not g31790 (n_15267, n16780);
  and g31791 (n16782, n_15266, n_15267);
  not g31792 (n_15268, n16781);
  not g31793 (n_15269, n16782);
  and g31794 (n16783, n_15268, n_15269);
  and g31795 (n16784, n16723, n16783);
  not g31796 (n_15270, n16723);
  not g31797 (n_15271, n16783);
  and g31798 (n16785, n_15270, n_15271);
  not g31799 (n_15272, n16784);
  not g31800 (n_15273, n16785);
  and g31801 (n16786, n_15272, n_15273);
  not g31802 (n_15274, n16660);
  and g31803 (n16787, n_15274, n16786);
  not g31804 (n_15275, n16786);
  and g31805 (n16788, n16660, n_15275);
  not g31806 (n_15276, n16787);
  not g31807 (n_15277, n16788);
  and g31808 (n16789, n_15276, n_15277);
  not g31809 (n_15278, n16659);
  not g31810 (n_15279, n16789);
  and g31811 (n16790, n_15278, n_15279);
  and g31812 (n16791, n16659, n16789);
  or g31813 (\asquared[98] , n16790, n16791);
  and g31814 (n16793, n_15269, n_15272);
  and g31815 (n16794, n_15258, n_15263);
  and g31816 (n16795, n_15195, n_15199);
  and g31817 (n16796, n_15155, n_15160);
  and g31818 (n16797, n16795, n16796);
  not g31819 (n_15280, n16795);
  not g31820 (n_15281, n16796);
  and g31821 (n16798, n_15280, n_15281);
  not g31822 (n_15282, n16797);
  not g31823 (n_15283, n16798);
  and g31824 (n16799, n_15282, n_15283);
  and g31825 (n16800, n_15238, n_15253);
  not g31826 (n_15284, n16799);
  and g31827 (n16801, n_15284, n16800);
  not g31828 (n_15285, n16800);
  and g31829 (n16802, n16799, n_15285);
  not g31830 (n_15286, n16801);
  not g31831 (n_15287, n16802);
  and g31832 (n16803, n_15286, n_15287);
  and g31833 (n16804, n16733, n16745);
  not g31834 (n_15288, n16733);
  not g31835 (n_15289, n16745);
  and g31836 (n16805, n_15288, n_15289);
  not g31837 (n_15290, n16804);
  not g31838 (n_15291, n16805);
  and g31839 (n16806, n_15290, n_15291);
  not g31840 (n_15292, n16806);
  and g31841 (n16807, n16764, n_15292);
  not g31842 (n_15293, n16764);
  and g31843 (n16808, n_15293, n16806);
  not g31844 (n_15294, n16807);
  not g31845 (n_15295, n16808);
  and g31846 (n16809, n_15294, n_15295);
  and g31847 (n16810, n_15185, n_15191);
  not g31848 (n_15296, n16809);
  and g31849 (n16811, n_15296, n16810);
  not g31850 (n_15297, n16810);
  and g31851 (n16812, n16809, n_15297);
  not g31852 (n_15298, n16811);
  not g31853 (n_15299, n16812);
  and g31854 (n16813, n_15298, n_15299);
  and g31855 (n16814, \a[39] , \a[59] );
  and g31856 (n16815, \a[40] , \a[58] );
  not g31857 (n_15300, n16814);
  not g31858 (n_15301, n16815);
  and g31859 (n16816, n_15300, n_15301);
  and g31860 (n16817, n4171, n8987);
  not g31861 (n_15302, n16817);
  not g31864 (n_15303, n16816);
  not g31866 (n_15304, n16820);
  and g31867 (n16821, n_15302, n_15304);
  and g31868 (n16822, n_15303, n16821);
  and g31869 (n16823, \a[53] , n_15304);
  and g31870 (n16824, \a[45] , n16823);
  not g31871 (n_15305, n16822);
  not g31872 (n_15306, n16824);
  and g31873 (n16825, n_15305, n_15306);
  and g31874 (n16826, n6252, n6564);
  and g31875 (n16827, n5666, n6968);
  and g31876 (n16828, \a[48] , \a[52] );
  and g31877 (n16829, n16557, n16828);
  not g31878 (n_15307, n16827);
  not g31879 (n_15308, n16829);
  and g31880 (n16830, n_15307, n_15308);
  not g31881 (n_15309, n16826);
  not g31882 (n_15310, n16830);
  and g31883 (n16831, n_15309, n_15310);
  not g31884 (n_15311, n16831);
  and g31885 (n16832, \a[52] , n_15311);
  and g31886 (n16833, \a[46] , n16832);
  and g31887 (n16834, n_15309, n_15311);
  not g31888 (n_15312, n5888);
  not g31889 (n_15313, n9127);
  and g31890 (n16835, n_15312, n_15313);
  not g31891 (n_15314, n16835);
  and g31892 (n16836, n16834, n_15314);
  not g31893 (n_15315, n16833);
  not g31894 (n_15316, n16836);
  and g31895 (n16837, n_15315, n_15316);
  not g31896 (n_15317, n16825);
  not g31897 (n_15318, n16837);
  and g31898 (n16838, n_15317, n_15318);
  not g31899 (n_15319, n16838);
  and g31900 (n16839, n_15317, n_15319);
  and g31901 (n16840, n_15318, n_15319);
  not g31902 (n_15320, n16839);
  not g31903 (n_15321, n16840);
  and g31904 (n16841, n_15320, n_15321);
  and g31905 (n16842, n3687, n9721);
  and g31906 (n16843, \a[37] , \a[61] );
  not g31907 (n_15322, n11588);
  not g31908 (n_15323, n16843);
  and g31909 (n16844, n_15322, n_15323);
  not g31910 (n_15324, n16842);
  not g31911 (n_15325, n16844);
  and g31912 (n16845, n_15324, n_15325);
  not g31913 (n_15326, n16680);
  and g31914 (n16846, n_15326, n16845);
  not g31915 (n_15327, n16845);
  and g31916 (n16847, n16680, n_15327);
  not g31917 (n_15328, n16846);
  not g31918 (n_15329, n16847);
  and g31919 (n16848, n_15328, n_15329);
  and g31920 (n16849, n16841, n16848);
  not g31921 (n_15330, n16841);
  not g31922 (n_15331, n16848);
  and g31923 (n16850, n_15330, n_15331);
  not g31924 (n_15332, n16849);
  not g31925 (n_15333, n16850);
  and g31926 (n16851, n_15332, n_15333);
  not g31927 (n_15334, n16851);
  and g31928 (n16852, n16813, n_15334);
  not g31929 (n_15335, n16852);
  and g31930 (n16853, n16813, n_15335);
  and g31931 (n16854, n_15334, n_15335);
  not g31932 (n_15336, n16853);
  not g31933 (n_15337, n16854);
  and g31934 (n16855, n_15336, n_15337);
  not g31935 (n_15338, n16855);
  and g31936 (n16856, n16803, n_15338);
  not g31937 (n_15339, n16803);
  and g31938 (n16857, n_15339, n16855);
  not g31939 (n_15340, n16794);
  not g31940 (n_15341, n16857);
  and g31941 (n16858, n_15340, n_15341);
  not g31942 (n_15342, n16856);
  and g31943 (n16859, n_15342, n16858);
  not g31944 (n_15343, n16859);
  and g31945 (n16860, n_15340, n_15343);
  and g31946 (n16861, n_15342, n_15343);
  and g31947 (n16862, n_15341, n16861);
  not g31948 (n_15344, n16860);
  not g31949 (n_15345, n16862);
  and g31950 (n16863, n_15344, n_15345);
  and g31951 (n16864, n_15210, n_15215);
  and g31952 (n16865, n_15203, n_15206);
  and g31953 (n16866, n5296, n7701);
  and g31954 (n16867, \a[43] , \a[55] );
  and g31955 (n16868, \a[44] , \a[54] );
  not g31956 (n_15346, n16867);
  not g31957 (n_15347, n16868);
  and g31958 (n16869, n_15346, n_15347);
  not g31959 (n_15348, n16866);
  not g31960 (n_15349, n16869);
  and g31961 (n16870, n_15348, n_15349);
  and g31962 (n16871, \a[35] , \a[63] );
  not g31963 (n_15350, n16870);
  not g31964 (n_15351, n16871);
  and g31965 (n16872, n_15350, n_15351);
  and g31966 (n16873, n16870, n16871);
  not g31967 (n_15352, n16872);
  not g31968 (n_15353, n16873);
  and g31969 (n16874, n_15352, n_15353);
  not g31970 (n_15354, n16694);
  and g31971 (n16875, n_15354, n16874);
  not g31972 (n_15355, n16874);
  and g31973 (n16876, n16694, n_15355);
  not g31974 (n_15356, n16875);
  not g31975 (n_15357, n16876);
  and g31976 (n16877, n_15356, n_15357);
  and g31977 (n16878, \a[38] , \a[60] );
  and g31978 (n16879, \a[41] , \a[57] );
  and g31979 (n16880, \a[42] , \a[56] );
  not g31980 (n_15358, n16879);
  not g31981 (n_15359, n16880);
  and g31982 (n16881, n_15358, n_15359);
  and g31983 (n16882, n5344, n8200);
  not g31984 (n_15360, n16882);
  and g31985 (n16883, n16878, n_15360);
  not g31986 (n_15361, n16881);
  and g31987 (n16884, n_15361, n16883);
  not g31988 (n_15362, n16884);
  and g31989 (n16885, n16878, n_15362);
  and g31990 (n16886, n_15360, n_15362);
  and g31991 (n16887, n_15361, n16886);
  not g31992 (n_15363, n16885);
  not g31993 (n_15364, n16887);
  and g31994 (n16888, n_15363, n_15364);
  not g31995 (n_15365, n16888);
  and g31996 (n16889, n16877, n_15365);
  not g31997 (n_15366, n16889);
  and g31998 (n16890, n16877, n_15366);
  and g31999 (n16891, n_15365, n_15366);
  not g32000 (n_15367, n16890);
  not g32001 (n_15368, n16891);
  and g32002 (n16892, n_15367, n_15368);
  and g32003 (n16893, n_15164, n_15167);
  not g32004 (n_15369, n16892);
  not g32005 (n_15370, n16893);
  and g32006 (n16894, n_15369, n_15370);
  not g32007 (n_15371, n16894);
  and g32008 (n16895, n_15369, n_15371);
  and g32009 (n16896, n_15370, n_15371);
  not g32010 (n_15372, n16895);
  not g32011 (n_15373, n16896);
  and g32012 (n16897, n_15372, n_15373);
  not g32013 (n_15374, n16865);
  not g32014 (n_15375, n16897);
  and g32015 (n16898, n_15374, n_15375);
  and g32016 (n16899, n16865, n_15373);
  and g32017 (n16900, n_15372, n16899);
  not g32018 (n_15376, n16898);
  not g32019 (n_15377, n16900);
  and g32020 (n16901, n_15376, n_15377);
  not g32021 (n_15378, n16864);
  and g32022 (n16902, n_15378, n16901);
  not g32023 (n_15379, n16902);
  and g32024 (n16903, n_15378, n_15379);
  and g32025 (n16904, n16901, n_15379);
  not g32026 (n_15380, n16903);
  not g32027 (n_15381, n16904);
  and g32028 (n16905, n_15380, n_15381);
  not g32029 (n_15382, n16863);
  not g32030 (n_15383, n16905);
  and g32031 (n16906, n_15382, n_15383);
  and g32032 (n16907, n16863, n_15381);
  and g32033 (n16908, n_15380, n16907);
  not g32034 (n_15384, n16906);
  not g32035 (n_15385, n16908);
  and g32036 (n16909, n_15384, n_15385);
  not g32037 (n_15386, n16909);
  and g32038 (n16910, n16793, n_15386);
  not g32039 (n_15387, n16793);
  and g32040 (n16911, n_15387, n16909);
  not g32041 (n_15388, n16910);
  not g32042 (n_15389, n16911);
  and g32043 (n16912, n_15388, n_15389);
  and g32044 (n16913, n_15278, n_15277);
  not g32045 (n_15390, n16913);
  and g32046 (n16914, n_15276, n_15390);
  not g32047 (n_15391, n16912);
  and g32048 (n16915, n_15391, n16914);
  not g32049 (n_15392, n16914);
  and g32050 (n16916, n16912, n_15392);
  not g32051 (n_15393, n16915);
  not g32052 (n_15394, n16916);
  and g32053 (\asquared[99] , n_15393, n_15394);
  and g32054 (n16918, n_15379, n_15384);
  and g32055 (n16919, n_15371, n_15376);
  and g32056 (n16920, n_15291, n_15295);
  and g32057 (n16921, \a[50] , \a[62] );
  and g32058 (n16922, \a[37] , n16921);
  not g32059 (n_15395, n16922);
  and g32060 (n16923, n6325, n_15395);
  not g32061 (n_15396, n16923);
  and g32062 (n16924, n6325, n_15396);
  and g32063 (n16925, n_15395, n_15396);
  and g32064 (n16926, \a[37] , \a[62] );
  not g32065 (n_15397, \a[50] );
  not g32066 (n_15398, n16926);
  and g32067 (n16927, n_15397, n_15398);
  not g32068 (n_15399, n16927);
  and g32069 (n16928, n16925, n_15399);
  not g32070 (n_15400, n16924);
  not g32071 (n_15401, n16928);
  and g32072 (n16929, n_15400, n_15401);
  not g32073 (n_15402, n16920);
  not g32074 (n_15403, n16929);
  and g32075 (n16930, n_15402, n_15403);
  not g32076 (n_15404, n16930);
  and g32077 (n16931, n_15402, n_15404);
  and g32078 (n16932, n_15403, n_15404);
  not g32079 (n_15405, n16931);
  not g32080 (n_15406, n16932);
  and g32081 (n16933, n_15405, n_15406);
  and g32082 (n16934, n_15356, n_15366);
  and g32083 (n16935, n16933, n16934);
  not g32084 (n_15407, n16933);
  not g32085 (n_15408, n16934);
  and g32086 (n16936, n_15407, n_15408);
  not g32087 (n_15409, n16935);
  not g32088 (n_15410, n16936);
  and g32089 (n16937, n_15409, n_15410);
  and g32090 (n16938, n_15324, n_15328);
  and g32091 (n16939, n16886, n16938);
  not g32092 (n_15411, n16886);
  not g32093 (n_15412, n16938);
  and g32094 (n16940, n_15411, n_15412);
  not g32095 (n_15413, n16939);
  not g32096 (n_15414, n16940);
  and g32097 (n16941, n_15413, n_15414);
  and g32098 (n16942, n5083, n9512);
  and g32099 (n16943, n8936, n11634);
  and g32100 (n16944, n3530, n9909);
  not g32101 (n_15415, n16943);
  not g32102 (n_15416, n16944);
  and g32103 (n16945, n_15415, n_15416);
  not g32104 (n_15417, n16942);
  not g32105 (n_15418, n16945);
  and g32106 (n16946, n_15417, n_15418);
  not g32107 (n_15419, n16946);
  and g32108 (n16947, \a[63] , n_15419);
  and g32109 (n16948, \a[36] , n16947);
  and g32110 (n16949, n_15417, n_15419);
  and g32111 (n16950, \a[38] , \a[61] );
  and g32112 (n16951, \a[39] , \a[60] );
  not g32113 (n_15420, n16950);
  not g32114 (n_15421, n16951);
  and g32115 (n16952, n_15420, n_15421);
  not g32116 (n_15422, n16952);
  and g32117 (n16953, n16949, n_15422);
  not g32118 (n_15423, n16948);
  not g32119 (n_15424, n16953);
  and g32120 (n16954, n_15423, n_15424);
  not g32121 (n_15425, n16954);
  and g32122 (n16955, n16941, n_15425);
  not g32123 (n_15426, n16955);
  and g32124 (n16956, n16941, n_15426);
  and g32125 (n16957, n_15425, n_15426);
  not g32126 (n_15427, n16956);
  not g32127 (n_15428, n16957);
  and g32128 (n16958, n_15427, n_15428);
  and g32129 (n16959, n16821, n16834);
  not g32130 (n_15429, n16821);
  not g32131 (n_15430, n16834);
  and g32132 (n16960, n_15429, n_15430);
  not g32133 (n_15431, n16959);
  not g32134 (n_15432, n16960);
  and g32135 (n16961, n_15431, n_15432);
  and g32136 (n16962, n_15348, n_15353);
  not g32137 (n_15433, n16961);
  and g32138 (n16963, n_15433, n16962);
  not g32139 (n_15434, n16962);
  and g32140 (n16964, n16961, n_15434);
  not g32141 (n_15435, n16963);
  not g32142 (n_15436, n16964);
  and g32143 (n16965, n_15435, n_15436);
  and g32144 (n16966, n_15330, n16848);
  not g32145 (n_15437, n16966);
  and g32146 (n16967, n_15319, n_15437);
  not g32147 (n_15438, n16967);
  and g32148 (n16968, n16965, n_15438);
  not g32149 (n_15439, n16965);
  and g32150 (n16969, n_15439, n16967);
  not g32151 (n_15440, n16968);
  not g32152 (n_15441, n16969);
  and g32153 (n16970, n_15440, n_15441);
  not g32154 (n_15442, n16958);
  not g32155 (n_15443, n16970);
  and g32156 (n16971, n_15442, n_15443);
  and g32157 (n16972, n16958, n16970);
  not g32158 (n_15444, n16971);
  not g32159 (n_15445, n16972);
  and g32160 (n16973, n_15444, n_15445);
  not g32161 (n_15446, n16973);
  and g32162 (n16974, n16937, n_15446);
  not g32163 (n_15447, n16937);
  and g32164 (n16975, n_15447, n16973);
  not g32165 (n_15448, n16974);
  not g32166 (n_15449, n16975);
  and g32167 (n16976, n_15448, n_15449);
  not g32168 (n_15450, n16919);
  and g32169 (n16977, n_15450, n16976);
  not g32170 (n_15451, n16976);
  and g32171 (n16978, n16919, n_15451);
  not g32172 (n_15452, n16977);
  not g32173 (n_15453, n16978);
  and g32174 (n16979, n_15452, n_15453);
  and g32175 (n16980, \a[41] , \a[58] );
  not g32176 (n_15454, n9490);
  not g32177 (n_15455, n16980);
  and g32178 (n16981, n_15454, n_15455);
  and g32179 (n16982, n5413, n8987);
  and g32180 (n16983, \a[44] , \a[59] );
  and g32181 (n16984, n16466, n16983);
  not g32182 (n_15456, n16982);
  not g32183 (n_15457, n16984);
  and g32184 (n16985, n_15456, n_15457);
  and g32185 (n16986, n9490, n16980);
  not g32186 (n_15458, n16985);
  not g32187 (n_15459, n16986);
  and g32188 (n16987, n_15458, n_15459);
  not g32189 (n_15460, n16987);
  and g32190 (n16988, n_15459, n_15460);
  not g32191 (n_15461, n16981);
  and g32192 (n16989, n_15461, n16988);
  and g32193 (n16990, \a[59] , n_15460);
  and g32194 (n16991, \a[40] , n16990);
  not g32195 (n_15462, n16989);
  not g32196 (n_15463, n16991);
  and g32197 (n16992, n_15462, n_15463);
  and g32198 (n16993, n5666, n7433);
  and g32199 (n16994, n5250, n10905);
  and g32200 (n16995, n5560, n7699);
  not g32201 (n_15464, n16994);
  not g32202 (n_15465, n16995);
  and g32203 (n16996, n_15464, n_15465);
  not g32204 (n_15466, n16993);
  not g32205 (n_15467, n16996);
  and g32206 (n16997, n_15466, n_15467);
  not g32207 (n_15468, n16997);
  and g32208 (n16998, \a[54] , n_15468);
  and g32209 (n16999, \a[45] , n16998);
  and g32210 (n17000, n_15466, n_15468);
  and g32211 (n17001, \a[46] , \a[53] );
  not g32212 (n_15469, n9428);
  not g32213 (n_15470, n17001);
  and g32214 (n17002, n_15469, n_15470);
  not g32215 (n_15471, n17002);
  and g32216 (n17003, n17000, n_15471);
  not g32217 (n_15472, n16999);
  not g32218 (n_15473, n17003);
  and g32219 (n17004, n_15472, n_15473);
  not g32220 (n_15474, n16992);
  not g32221 (n_15475, n17004);
  and g32222 (n17005, n_15474, n_15475);
  not g32223 (n_15476, n17005);
  and g32224 (n17006, n_15474, n_15476);
  and g32225 (n17007, n_15475, n_15476);
  not g32226 (n_15477, n17006);
  not g32227 (n_15478, n17007);
  and g32228 (n17008, n_15477, n_15478);
  and g32229 (n17009, \a[48] , \a[51] );
  and g32230 (n17010, \a[42] , \a[57] );
  and g32231 (n17011, \a[43] , \a[56] );
  not g32232 (n_15479, n17010);
  not g32233 (n_15480, n17011);
  and g32234 (n17012, n_15479, n_15480);
  and g32235 (n17013, n5018, n8200);
  not g32236 (n_15481, n17013);
  and g32237 (n17014, n17009, n_15481);
  not g32238 (n_15482, n17012);
  and g32239 (n17015, n_15482, n17014);
  not g32240 (n_15483, n17015);
  and g32241 (n17016, n17009, n_15483);
  and g32242 (n17017, n_15481, n_15483);
  and g32243 (n17018, n_15482, n17017);
  not g32244 (n_15484, n17016);
  not g32245 (n_15485, n17018);
  and g32246 (n17019, n_15484, n_15485);
  not g32247 (n_15486, n17008);
  not g32248 (n_15487, n17019);
  and g32249 (n17020, n_15486, n_15487);
  not g32250 (n_15488, n17020);
  and g32251 (n17021, n_15486, n_15488);
  and g32252 (n17022, n_15487, n_15488);
  not g32253 (n_15489, n17021);
  not g32254 (n_15490, n17022);
  and g32255 (n17023, n_15489, n_15490);
  and g32256 (n17024, n_15283, n_15287);
  and g32257 (n17025, n17023, n17024);
  not g32258 (n_15491, n17023);
  not g32259 (n_15492, n17024);
  and g32260 (n17026, n_15491, n_15492);
  not g32261 (n_15493, n17025);
  not g32262 (n_15494, n17026);
  and g32263 (n17027, n_15493, n_15494);
  and g32264 (n17028, n_15299, n_15335);
  not g32265 (n_15495, n17027);
  and g32266 (n17029, n_15495, n17028);
  not g32267 (n_15496, n17028);
  and g32268 (n17030, n17027, n_15496);
  not g32269 (n_15497, n17029);
  not g32270 (n_15498, n17030);
  and g32271 (n17031, n_15497, n_15498);
  not g32272 (n_15499, n16861);
  and g32273 (n17032, n_15499, n17031);
  not g32274 (n_15500, n17032);
  and g32275 (n17033, n17031, n_15500);
  and g32276 (n17034, n_15499, n_15500);
  not g32277 (n_15501, n17033);
  not g32278 (n_15502, n17034);
  and g32279 (n17035, n_15501, n_15502);
  not g32280 (n_15503, n17035);
  and g32281 (n17036, n16979, n_15503);
  not g32282 (n_15504, n16979);
  and g32283 (n17037, n_15504, n_15502);
  and g32284 (n17038, n_15501, n17037);
  not g32285 (n_15505, n17036);
  not g32286 (n_15506, n17038);
  and g32287 (n17039, n_15505, n_15506);
  not g32288 (n_15507, n16918);
  and g32289 (n17040, n_15507, n17039);
  not g32290 (n_15508, n17039);
  and g32291 (n17041, n16918, n_15508);
  not g32292 (n_15509, n17040);
  not g32293 (n_15510, n17041);
  and g32294 (n17042, n_15509, n_15510);
  and g32295 (n17043, n_15388, n_15392);
  not g32296 (n_15511, n17043);
  and g32297 (n17044, n_15389, n_15511);
  not g32298 (n_15512, n17042);
  and g32299 (n17045, n_15512, n17044);
  not g32300 (n_15513, n17044);
  and g32301 (n17046, n17042, n_15513);
  not g32302 (n_15514, n17045);
  not g32303 (n_15515, n17046);
  and g32304 (\asquared[100] , n_15514, n_15515);
  and g32305 (n17048, n_15510, n_15513);
  not g32306 (n_15516, n17048);
  and g32307 (n17049, n_15509, n_15516);
  and g32308 (n17050, n_15500, n_15505);
  and g32309 (n17051, n_15432, n_15436);
  and g32310 (n17052, n6256, n6968);
  and g32311 (n17053, n6254, n7232);
  and g32312 (n17054, n6252, n7433);
  not g32313 (n_15517, n17053);
  not g32314 (n_15518, n17054);
  and g32315 (n17055, n_15517, n_15518);
  not g32316 (n_15519, n17052);
  not g32317 (n_15520, n17055);
  and g32318 (n17056, n_15519, n_15520);
  not g32319 (n_15521, n17056);
  and g32320 (n17057, \a[53] , n_15521);
  and g32321 (n17058, \a[47] , n17057);
  and g32322 (n17059, n_15519, n_15521);
  not g32323 (n_15522, n9934);
  not g32324 (n_15523, n16828);
  and g32325 (n17060, n_15522, n_15523);
  not g32326 (n_15524, n17060);
  and g32327 (n17061, n17059, n_15524);
  not g32328 (n_15525, n17058);
  not g32329 (n_15526, n17061);
  and g32330 (n17062, n_15525, n_15526);
  not g32331 (n_15527, n17051);
  not g32332 (n_15528, n17062);
  and g32333 (n17063, n_15527, n_15528);
  not g32334 (n_15529, n17063);
  and g32335 (n17064, n_15527, n_15529);
  and g32336 (n17065, n_15528, n_15529);
  not g32337 (n_15530, n17064);
  not g32338 (n_15531, n17065);
  and g32339 (n17066, n_15530, n_15531);
  and g32340 (n17067, n_15414, n_15426);
  and g32341 (n17068, n17066, n17067);
  not g32342 (n_15532, n17066);
  not g32343 (n_15533, n17067);
  and g32344 (n17069, n_15532, n_15533);
  not g32345 (n_15534, n17068);
  not g32346 (n_15535, n17069);
  and g32347 (n17070, n_15534, n_15535);
  and g32348 (n17071, n_15494, n_15498);
  not g32349 (n_15536, n17070);
  and g32350 (n17072, n_15536, n17071);
  not g32351 (n_15537, n17071);
  and g32352 (n17073, n17070, n_15537);
  not g32353 (n_15538, n17072);
  not g32354 (n_15539, n17073);
  and g32355 (n17074, n_15538, n_15539);
  and g32356 (n17075, n16949, n17000);
  not g32357 (n_15540, n16949);
  not g32358 (n_15541, n17000);
  and g32359 (n17076, n_15540, n_15541);
  not g32360 (n_15542, n17075);
  not g32361 (n_15543, n17076);
  and g32362 (n17077, n_15542, n_15543);
  not g32363 (n_15544, n17077);
  and g32364 (n17078, n16988, n_15544);
  not g32365 (n_15545, n16988);
  and g32366 (n17079, n_15545, n17077);
  not g32367 (n_15546, n17078);
  not g32368 (n_15547, n17079);
  and g32369 (n17080, n_15546, n_15547);
  and g32370 (n17081, n_15476, n_15488);
  not g32371 (n_15548, n17080);
  and g32372 (n17082, n_15548, n17081);
  not g32373 (n_15549, n17081);
  and g32374 (n17083, n17080, n_15549);
  not g32375 (n_15550, n17082);
  not g32376 (n_15551, n17083);
  and g32377 (n17084, n_15550, n_15551);
  and g32378 (n17085, \a[37] , \a[63] );
  not g32379 (n_15552, n16925);
  and g32380 (n17086, n_15552, n17085);
  not g32381 (n_15553, n17085);
  and g32382 (n17087, n16925, n_15553);
  not g32383 (n_15554, n17086);
  not g32384 (n_15555, n17087);
  and g32385 (n17088, n_15554, n_15555);
  not g32386 (n_15556, n17088);
  and g32387 (n17089, n17017, n_15556);
  not g32388 (n_15557, n17017);
  and g32389 (n17090, n_15557, n17088);
  not g32390 (n_15558, n17089);
  not g32391 (n_15559, n17090);
  and g32392 (n17091, n_15558, n_15559);
  and g32393 (n17092, n17084, n17091);
  not g32394 (n_15560, n17084);
  not g32395 (n_15561, n17091);
  and g32396 (n17093, n_15560, n_15561);
  not g32397 (n_15562, n17092);
  not g32398 (n_15563, n17093);
  and g32399 (n17094, n_15562, n_15563);
  and g32400 (n17095, n17074, n17094);
  not g32401 (n_15564, n17074);
  not g32402 (n_15565, n17094);
  and g32403 (n17096, n_15564, n_15565);
  not g32404 (n_15566, n17095);
  not g32405 (n_15567, n17096);
  and g32406 (n17097, n_15566, n_15567);
  and g32407 (n17098, n_15448, n_15452);
  and g32408 (n17099, n4171, n9512);
  and g32409 (n17100, n13544, n16878);
  and g32410 (n17101, n5083, n9721);
  not g32411 (n_15568, n17100);
  not g32412 (n_15569, n17101);
  and g32413 (n17102, n_15568, n_15569);
  not g32414 (n_15570, n17099);
  not g32415 (n_15571, n17102);
  and g32416 (n17103, n_15570, n_15571);
  not g32417 (n_15572, n17103);
  and g32418 (n17104, n_15570, n_15572);
  and g32419 (n17105, \a[39] , \a[61] );
  not g32420 (n_15573, n16523);
  not g32421 (n_15574, n17105);
  and g32422 (n17106, n_15573, n_15574);
  not g32423 (n_15575, n17106);
  and g32424 (n17107, n17104, n_15575);
  and g32425 (n17108, n12571, n_15572);
  not g32426 (n_15576, n17107);
  not g32427 (n_15577, n17108);
  and g32428 (n17109, n_15576, n_15577);
  and g32429 (n17110, n5713, n9161);
  and g32430 (n17111, n4811, n11718);
  and g32431 (n17112, n5296, n8200);
  not g32432 (n_15578, n17111);
  not g32433 (n_15579, n17112);
  and g32434 (n17113, n_15578, n_15579);
  not g32435 (n_15580, n17110);
  not g32436 (n_15581, n17113);
  and g32437 (n17114, n_15580, n_15581);
  not g32438 (n_15582, n17114);
  and g32439 (n17115, n10303, n_15582);
  not g32440 (n_15583, n9493);
  not g32441 (n_15584, n16167);
  and g32442 (n17116, n_15583, n_15584);
  and g32443 (n17117, n_15580, n_15582);
  not g32444 (n_15585, n17116);
  and g32445 (n17118, n_15585, n17117);
  not g32446 (n_15586, n17115);
  not g32447 (n_15587, n17118);
  and g32448 (n17119, n_15586, n_15587);
  not g32449 (n_15588, n17109);
  not g32450 (n_15589, n17119);
  and g32451 (n17120, n_15588, n_15589);
  not g32452 (n_15590, n17120);
  and g32453 (n17121, n_15588, n_15590);
  and g32454 (n17122, n_15589, n_15590);
  not g32455 (n_15591, n17121);
  not g32456 (n_15592, n17122);
  and g32457 (n17123, n_15591, n_15592);
  and g32458 (n17124, \a[41] , \a[59] );
  and g32459 (n17125, \a[42] , \a[58] );
  not g32460 (n_15593, n17124);
  not g32461 (n_15594, n17125);
  and g32462 (n17126, n_15593, n_15594);
  and g32463 (n17127, n5344, n8987);
  not g32464 (n_15595, n17127);
  and g32465 (n17128, n9414, n_15595);
  not g32466 (n_15596, n17126);
  and g32467 (n17129, n_15596, n17128);
  not g32468 (n_15597, n17129);
  and g32469 (n17130, n9414, n_15597);
  and g32470 (n17131, n_15595, n_15597);
  and g32471 (n17132, n_15596, n17131);
  not g32472 (n_15598, n17130);
  not g32473 (n_15599, n17132);
  and g32474 (n17133, n_15598, n_15599);
  not g32475 (n_15600, n17123);
  not g32476 (n_15601, n17133);
  and g32477 (n17134, n_15600, n_15601);
  not g32478 (n_15602, n17134);
  and g32479 (n17135, n_15600, n_15602);
  and g32480 (n17136, n_15601, n_15602);
  not g32481 (n_15603, n17135);
  not g32482 (n_15604, n17136);
  and g32483 (n17137, n_15603, n_15604);
  and g32484 (n17138, n_15404, n_15410);
  and g32485 (n17139, n17137, n17138);
  not g32486 (n_15605, n17137);
  not g32487 (n_15606, n17138);
  and g32488 (n17140, n_15605, n_15606);
  not g32489 (n_15607, n17139);
  not g32490 (n_15608, n17140);
  and g32491 (n17141, n_15607, n_15608);
  and g32492 (n17142, n_15442, n16970);
  not g32493 (n_15609, n17142);
  and g32494 (n17143, n_15440, n_15609);
  not g32495 (n_15610, n17143);
  and g32496 (n17144, n17141, n_15610);
  not g32497 (n_15611, n17141);
  and g32498 (n17145, n_15611, n17143);
  not g32499 (n_15612, n17144);
  not g32500 (n_15613, n17145);
  and g32501 (n17146, n_15612, n_15613);
  not g32502 (n_15614, n17098);
  and g32503 (n17147, n_15614, n17146);
  not g32504 (n_15615, n17146);
  and g32505 (n17148, n17098, n_15615);
  not g32506 (n_15616, n17147);
  not g32507 (n_15617, n17148);
  and g32508 (n17149, n_15616, n_15617);
  and g32509 (n17150, n17097, n17149);
  not g32510 (n_15618, n17097);
  not g32511 (n_15619, n17149);
  and g32512 (n17151, n_15618, n_15619);
  not g32513 (n_15620, n17150);
  not g32514 (n_15621, n17151);
  and g32515 (n17152, n_15620, n_15621);
  not g32516 (n_15622, n17050);
  and g32517 (n17153, n_15622, n17152);
  not g32518 (n_15623, n17152);
  and g32519 (n17154, n17050, n_15623);
  not g32520 (n_15624, n17153);
  not g32521 (n_15625, n17154);
  and g32522 (n17155, n_15624, n_15625);
  not g32523 (n_15626, n17155);
  and g32524 (n17156, n17049, n_15626);
  not g32525 (n_15627, n17049);
  and g32526 (n17157, n_15627, n_15625);
  and g32527 (n17158, n_15624, n17157);
  not g32528 (n_15628, n17156);
  not g32529 (n_15629, n17158);
  and g32530 (\asquared[101] , n_15628, n_15629);
  not g32531 (n_15630, n17157);
  and g32532 (n17160, n_15624, n_15630);
  and g32533 (n17161, n_15616, n_15620);
  and g32534 (n17162, n_15539, n_15566);
  and g32535 (n17163, \a[46] , \a[55] );
  and g32536 (n17164, \a[47] , \a[54] );
  not g32537 (n_15631, n17163);
  not g32538 (n_15632, n17164);
  and g32539 (n17165, n_15631, n_15632);
  and g32540 (n17166, n5666, n7701);
  not g32541 (n_15633, n17166);
  not g32544 (n_15634, n17165);
  not g32546 (n_15635, n17169);
  and g32547 (n17170, n_15633, n_15635);
  and g32548 (n17171, n_15634, n17170);
  and g32549 (n17172, \a[63] , n_15635);
  and g32550 (n17173, \a[38] , n17172);
  not g32551 (n_15636, n17171);
  not g32552 (n_15637, n17173);
  and g32553 (n17174, n_15636, n_15637);
  and g32554 (n17175, n4811, n7942);
  and g32555 (n17176, n13870, n15167);
  and g32556 (n17177, n5018, n8987);
  not g32557 (n_15638, n17176);
  not g32558 (n_15639, n17177);
  and g32559 (n17178, n_15638, n_15639);
  not g32560 (n_15640, n17175);
  not g32561 (n_15641, n17178);
  and g32562 (n17179, n_15640, n_15641);
  not g32563 (n_15642, n17179);
  and g32564 (n17180, \a[59] , n_15642);
  and g32565 (n17181, \a[42] , n17180);
  and g32566 (n17182, n_15640, n_15642);
  and g32567 (n17183, \a[43] , \a[58] );
  and g32568 (n17184, \a[45] , \a[56] );
  not g32569 (n_15643, n17183);
  not g32570 (n_15644, n17184);
  and g32571 (n17185, n_15643, n_15644);
  not g32572 (n_15645, n17185);
  and g32573 (n17186, n17182, n_15645);
  not g32574 (n_15646, n17181);
  not g32575 (n_15647, n17186);
  and g32576 (n17187, n_15646, n_15647);
  not g32577 (n_15648, n17174);
  not g32578 (n_15649, n17187);
  and g32579 (n17188, n_15648, n_15649);
  not g32580 (n_15650, n17188);
  and g32581 (n17189, n_15648, n_15650);
  and g32582 (n17190, n_15649, n_15650);
  not g32583 (n_15651, n17189);
  not g32584 (n_15652, n17190);
  and g32585 (n17191, n_15651, n_15652);
  and g32586 (n17192, n8700, n12601);
  and g32587 (n17193, n6256, n7433);
  and g32588 (n17194, \a[44] , \a[57] );
  and g32589 (n17195, n10439, n17194);
  not g32590 (n_15653, n17193);
  not g32591 (n_15654, n17195);
  and g32592 (n17196, n_15653, n_15654);
  not g32593 (n_15655, n17192);
  not g32594 (n_15656, n17196);
  and g32595 (n17197, n_15655, n_15656);
  not g32596 (n_15657, n17197);
  and g32597 (n17198, n10439, n_15657);
  and g32598 (n17199, n_15655, n_15657);
  and g32599 (n17200, \a[49] , \a[52] );
  not g32600 (n_15658, n17194);
  not g32601 (n_15659, n17200);
  and g32602 (n17201, n_15658, n_15659);
  not g32603 (n_15660, n17201);
  and g32604 (n17202, n17199, n_15660);
  not g32605 (n_15661, n17198);
  not g32606 (n_15662, n17202);
  and g32607 (n17203, n_15661, n_15662);
  not g32608 (n_15663, n17191);
  not g32609 (n_15664, n17203);
  and g32610 (n17204, n_15663, n_15664);
  not g32611 (n_15665, n17204);
  and g32612 (n17205, n_15663, n_15665);
  and g32613 (n17206, n_15664, n_15665);
  not g32614 (n_15666, n17205);
  not g32615 (n_15667, n17206);
  and g32616 (n17207, n_15666, n_15667);
  and g32617 (n17208, n_15529, n_15535);
  and g32618 (n17209, n17207, n17208);
  not g32619 (n_15668, n17207);
  not g32620 (n_15669, n17208);
  and g32621 (n17210, n_15668, n_15669);
  not g32622 (n_15670, n17209);
  not g32623 (n_15671, n17210);
  and g32624 (n17211, n_15670, n_15671);
  and g32625 (n17212, n_15554, n_15559);
  and g32626 (n17213, n5413, n9512);
  not g32627 (n_15672, n17213);
  and g32628 (n17214, \a[60] , n_15672);
  and g32629 (n17215, \a[41] , n17214);
  and g32630 (n17216, \a[61] , n_15672);
  and g32631 (n17217, \a[40] , n17216);
  not g32632 (n_15673, n17215);
  not g32633 (n_15674, n17217);
  and g32634 (n17218, n_15673, n_15674);
  not g32635 (n_15675, n17059);
  not g32636 (n_15676, n17218);
  and g32637 (n17219, n_15675, n_15676);
  not g32638 (n_15677, n17219);
  and g32639 (n17220, n_15675, n_15677);
  and g32640 (n17221, n_15676, n_15677);
  not g32641 (n_15678, n17220);
  not g32642 (n_15679, n17221);
  and g32643 (n17222, n_15678, n_15679);
  and g32644 (n17223, \a[62] , n7774);
  not g32645 (n_15680, n17223);
  and g32646 (n17224, n6564, n_15680);
  not g32647 (n_15681, n17224);
  and g32648 (n17225, n_15680, n_15681);
  and g32649 (n17226, \a[39] , \a[62] );
  not g32650 (n_15682, \a[51] );
  not g32651 (n_15683, n17226);
  and g32652 (n17227, n_15682, n_15683);
  not g32653 (n_15684, n17227);
  and g32654 (n17228, n17225, n_15684);
  and g32655 (n17229, n6564, n_15681);
  not g32656 (n_15685, n17228);
  not g32657 (n_15686, n17229);
  and g32658 (n17230, n_15685, n_15686);
  not g32659 (n_15687, n17222);
  not g32660 (n_15688, n17230);
  and g32661 (n17231, n_15687, n_15688);
  not g32662 (n_15689, n17231);
  and g32663 (n17232, n_15687, n_15689);
  and g32664 (n17233, n_15688, n_15689);
  not g32665 (n_15690, n17232);
  not g32666 (n_15691, n17233);
  and g32667 (n17234, n_15690, n_15691);
  not g32668 (n_15692, n17212);
  not g32669 (n_15693, n17234);
  and g32670 (n17235, n_15692, n_15693);
  not g32671 (n_15694, n17235);
  and g32672 (n17236, n_15692, n_15694);
  and g32673 (n17237, n_15693, n_15694);
  not g32674 (n_15695, n17236);
  not g32675 (n_15696, n17237);
  and g32676 (n17238, n_15695, n_15696);
  not g32677 (n_15697, n17238);
  and g32678 (n17239, n17211, n_15697);
  not g32679 (n_15698, n17211);
  and g32680 (n17240, n_15698, n17238);
  not g32681 (n_15699, n17162);
  not g32682 (n_15700, n17240);
  and g32683 (n17241, n_15699, n_15700);
  not g32684 (n_15701, n17239);
  and g32685 (n17242, n_15701, n17241);
  not g32686 (n_15702, n17242);
  and g32687 (n17243, n_15699, n_15702);
  and g32688 (n17244, n_15700, n_15702);
  and g32689 (n17245, n_15701, n17244);
  not g32690 (n_15703, n17243);
  not g32691 (n_15704, n17245);
  and g32692 (n17246, n_15703, n_15704);
  and g32693 (n17247, n_15608, n_15612);
  and g32694 (n17248, n_15551, n_15562);
  not g32695 (n_15705, n17247);
  not g32696 (n_15706, n17248);
  and g32697 (n17249, n_15705, n_15706);
  not g32698 (n_15707, n17249);
  and g32699 (n17250, n_15705, n_15707);
  and g32700 (n17251, n_15706, n_15707);
  not g32701 (n_15708, n17250);
  not g32702 (n_15709, n17251);
  and g32703 (n17252, n_15708, n_15709);
  and g32704 (n17253, n17104, n17131);
  not g32705 (n_15710, n17104);
  not g32706 (n_15711, n17131);
  and g32707 (n17254, n_15710, n_15711);
  not g32708 (n_15712, n17253);
  not g32709 (n_15713, n17254);
  and g32710 (n17255, n_15712, n_15713);
  not g32711 (n_15714, n17255);
  and g32712 (n17256, n17117, n_15714);
  not g32713 (n_15715, n17117);
  and g32714 (n17257, n_15715, n17255);
  not g32715 (n_15716, n17256);
  not g32716 (n_15717, n17257);
  and g32717 (n17258, n_15716, n_15717);
  and g32718 (n17259, n_15590, n_15602);
  and g32719 (n17260, n_15543, n_15547);
  and g32720 (n17261, n17259, n17260);
  not g32721 (n_15718, n17259);
  not g32722 (n_15719, n17260);
  and g32723 (n17262, n_15718, n_15719);
  not g32724 (n_15720, n17261);
  not g32725 (n_15721, n17262);
  and g32726 (n17263, n_15720, n_15721);
  and g32727 (n17264, n17258, n17263);
  not g32728 (n_15722, n17258);
  not g32729 (n_15723, n17263);
  and g32730 (n17265, n_15722, n_15723);
  not g32731 (n_15724, n17264);
  not g32732 (n_15725, n17265);
  and g32733 (n17266, n_15724, n_15725);
  not g32734 (n_15726, n17252);
  and g32735 (n17267, n_15726, n17266);
  not g32736 (n_15727, n17267);
  and g32737 (n17268, n_15726, n_15727);
  and g32738 (n17269, n17266, n_15727);
  not g32739 (n_15728, n17268);
  not g32740 (n_15729, n17269);
  and g32741 (n17270, n_15728, n_15729);
  not g32742 (n_15730, n17246);
  and g32743 (n17271, n_15730, n17270);
  not g32744 (n_15731, n17270);
  and g32745 (n17272, n17246, n_15731);
  not g32746 (n_15732, n17271);
  not g32747 (n_15733, n17272);
  and g32748 (n17273, n_15732, n_15733);
  not g32749 (n_15734, n17161);
  not g32750 (n_15735, n17273);
  and g32751 (n17274, n_15734, n_15735);
  and g32752 (n17275, n17161, n17273);
  not g32753 (n_15736, n17274);
  not g32754 (n_15737, n17275);
  and g32755 (n17276, n_15736, n_15737);
  not g32756 (n_15738, n17160);
  not g32757 (n_15739, n17276);
  and g32758 (n17277, n_15738, n_15739);
  and g32759 (n17278, n17160, n17276);
  or g32760 (\asquared[102] , n17277, n17278);
  and g32761 (n17280, n_15738, n_15737);
  not g32762 (n_15740, n17280);
  and g32763 (n17281, n_15736, n_15740);
  and g32764 (n17282, n_15730, n_15731);
  not g32765 (n_15741, n17282);
  and g32766 (n17283, n_15702, n_15741);
  and g32767 (n17284, n_15707, n_15727);
  and g32768 (n17285, n_15672, n_15677);
  and g32769 (n17286, n17182, n17285);
  not g32770 (n_15742, n17182);
  not g32771 (n_15743, n17285);
  and g32772 (n17287, n_15742, n_15743);
  not g32773 (n_15744, n17286);
  not g32774 (n_15745, n17287);
  and g32775 (n17288, n_15744, n_15745);
  and g32776 (n17289, n5344, n9512);
  and g32777 (n17290, n11634, n13971);
  and g32778 (n17291, n3984, n9909);
  not g32779 (n_15746, n17290);
  not g32780 (n_15747, n17291);
  and g32781 (n17292, n_15746, n_15747);
  not g32782 (n_15748, n17289);
  not g32783 (n_15749, n17292);
  and g32784 (n17293, n_15748, n_15749);
  not g32785 (n_15750, n17293);
  and g32786 (n17294, \a[63] , n_15750);
  and g32787 (n17295, \a[39] , n17294);
  and g32788 (n17296, n_15748, n_15750);
  and g32789 (n17297, \a[41] , \a[61] );
  and g32790 (n17298, \a[42] , \a[60] );
  not g32791 (n_15751, n17297);
  not g32792 (n_15752, n17298);
  and g32793 (n17299, n_15751, n_15752);
  not g32794 (n_15753, n17299);
  and g32795 (n17300, n17296, n_15753);
  not g32796 (n_15754, n17295);
  not g32797 (n_15755, n17300);
  and g32798 (n17301, n_15754, n_15755);
  not g32799 (n_15756, n17301);
  and g32800 (n17302, n17288, n_15756);
  not g32801 (n_15757, n17302);
  and g32802 (n17303, n17288, n_15757);
  and g32803 (n17304, n_15756, n_15757);
  not g32804 (n_15758, n17303);
  not g32805 (n_15759, n17304);
  and g32806 (n17305, n_15758, n_15759);
  and g32807 (n17306, n_15689, n_15694);
  and g32808 (n17307, n17305, n17306);
  not g32809 (n_15760, n17305);
  not g32810 (n_15761, n17306);
  and g32811 (n17308, n_15760, n_15761);
  not g32812 (n_15762, n17307);
  not g32813 (n_15763, n17308);
  and g32814 (n17309, n_15762, n_15763);
  and g32815 (n17310, \a[43] , \a[59] );
  and g32816 (n17311, \a[44] , \a[58] );
  not g32817 (n_15764, n17310);
  not g32818 (n_15765, n17311);
  and g32819 (n17312, n_15764, n_15765);
  and g32820 (n17313, n5296, n8987);
  not g32821 (n_15766, n17313);
  and g32822 (n17314, n13544, n_15766);
  not g32823 (n_15767, n17312);
  and g32824 (n17315, n_15767, n17314);
  not g32825 (n_15768, n17315);
  and g32826 (n17316, n_15766, n_15768);
  and g32827 (n17317, n_15767, n17316);
  and g32828 (n17318, n13544, n_15768);
  not g32829 (n_15769, n17317);
  not g32830 (n_15770, n17318);
  and g32831 (n17319, n_15769, n_15770);
  and g32832 (n17320, n5666, n9161);
  and g32833 (n17321, n5250, n11718);
  and g32834 (n17322, n5560, n8200);
  not g32835 (n_15771, n17321);
  not g32836 (n_15772, n17322);
  and g32837 (n17323, n_15771, n_15772);
  not g32838 (n_15773, n17320);
  not g32839 (n_15774, n17323);
  and g32840 (n17324, n_15773, n_15774);
  not g32841 (n_15775, n17324);
  and g32842 (n17325, \a[57] , n_15775);
  and g32843 (n17326, \a[45] , n17325);
  and g32844 (n17327, \a[46] , \a[56] );
  and g32845 (n17328, \a[47] , \a[55] );
  not g32846 (n_15776, n17327);
  not g32847 (n_15777, n17328);
  and g32848 (n17329, n_15776, n_15777);
  and g32849 (n17330, n_15773, n_15775);
  not g32850 (n_15778, n17329);
  and g32851 (n17331, n_15778, n17330);
  not g32852 (n_15779, n17326);
  not g32853 (n_15780, n17331);
  and g32854 (n17332, n_15779, n_15780);
  not g32855 (n_15781, n17319);
  not g32856 (n_15782, n17332);
  and g32857 (n17333, n_15781, n_15782);
  not g32858 (n_15783, n17333);
  and g32859 (n17334, n_15781, n_15783);
  and g32860 (n17335, n_15782, n_15783);
  not g32861 (n_15784, n17334);
  not g32862 (n_15785, n17335);
  and g32863 (n17336, n_15784, n_15785);
  and g32864 (n17337, n6325, n7433);
  and g32865 (n17338, n5888, n10905);
  and g32866 (n17339, n6256, n7699);
  not g32867 (n_15786, n17338);
  not g32868 (n_15787, n17339);
  and g32869 (n17340, n_15786, n_15787);
  not g32870 (n_15788, n17337);
  not g32871 (n_15789, n17340);
  and g32872 (n17341, n_15788, n_15789);
  not g32873 (n_15790, n17341);
  and g32874 (n17342, \a[54] , n_15790);
  and g32875 (n17343, \a[48] , n17342);
  and g32876 (n17344, n_15788, n_15790);
  and g32877 (n17345, \a[49] , \a[53] );
  not g32878 (n_15791, n6966);
  not g32879 (n_15792, n17345);
  and g32880 (n17346, n_15791, n_15792);
  not g32881 (n_15793, n17346);
  and g32882 (n17347, n17344, n_15793);
  not g32883 (n_15794, n17343);
  not g32884 (n_15795, n17347);
  and g32885 (n17348, n_15794, n_15795);
  not g32886 (n_15796, n17336);
  not g32887 (n_15797, n17348);
  and g32888 (n17349, n_15796, n_15797);
  not g32889 (n_15798, n17349);
  and g32890 (n17350, n_15796, n_15798);
  and g32891 (n17351, n_15797, n_15798);
  not g32892 (n_15799, n17350);
  not g32893 (n_15800, n17351);
  and g32894 (n17352, n_15799, n_15800);
  not g32895 (n_15801, n17352);
  and g32896 (n17353, n17309, n_15801);
  not g32897 (n_15802, n17309);
  and g32898 (n17354, n_15802, n17352);
  not g32899 (n_15803, n17284);
  not g32900 (n_15804, n17354);
  and g32901 (n17355, n_15803, n_15804);
  not g32902 (n_15805, n17353);
  and g32903 (n17356, n_15805, n17355);
  not g32904 (n_15806, n17356);
  and g32905 (n17357, n_15803, n_15806);
  and g32906 (n17358, n_15804, n_15806);
  and g32907 (n17359, n_15805, n17358);
  not g32908 (n_15807, n17357);
  not g32909 (n_15808, n17359);
  and g32910 (n17360, n_15807, n_15808);
  and g32911 (n17361, n17199, n17225);
  not g32912 (n_15809, n17199);
  not g32913 (n_15810, n17225);
  and g32914 (n17362, n_15809, n_15810);
  not g32915 (n_15811, n17361);
  not g32916 (n_15812, n17362);
  and g32917 (n17363, n_15811, n_15812);
  not g32918 (n_15813, n17363);
  and g32919 (n17364, n17170, n_15813);
  not g32920 (n_15814, n17170);
  and g32921 (n17365, n_15814, n17363);
  not g32922 (n_15815, n17364);
  not g32923 (n_15816, n17365);
  and g32924 (n17366, n_15815, n_15816);
  and g32925 (n17367, n_15713, n_15717);
  not g32926 (n_15817, n17366);
  and g32927 (n17368, n_15817, n17367);
  not g32928 (n_15818, n17367);
  and g32929 (n17369, n17366, n_15818);
  not g32930 (n_15819, n17368);
  not g32931 (n_15820, n17369);
  and g32932 (n17370, n_15819, n_15820);
  and g32933 (n17371, n_15650, n_15665);
  not g32934 (n_15821, n17370);
  and g32935 (n17372, n_15821, n17371);
  not g32936 (n_15822, n17371);
  and g32937 (n17373, n17370, n_15822);
  not g32938 (n_15823, n17372);
  not g32939 (n_15824, n17373);
  and g32940 (n17374, n_15823, n_15824);
  and g32941 (n17375, n_15671, n_15701);
  and g32942 (n17376, n_15721, n_15724);
  not g32943 (n_15825, n17375);
  not g32944 (n_15826, n17376);
  and g32945 (n17377, n_15825, n_15826);
  not g32946 (n_15827, n17377);
  and g32947 (n17378, n_15825, n_15827);
  and g32948 (n17379, n_15826, n_15827);
  not g32949 (n_15828, n17378);
  not g32950 (n_15829, n17379);
  and g32951 (n17380, n_15828, n_15829);
  not g32952 (n_15830, n17380);
  and g32953 (n17381, n17374, n_15830);
  not g32954 (n_15831, n17374);
  and g32955 (n17382, n_15831, n17380);
  not g32956 (n_15832, n17360);
  not g32957 (n_15833, n17382);
  and g32958 (n17383, n_15832, n_15833);
  not g32959 (n_15834, n17381);
  and g32960 (n17384, n_15834, n17383);
  not g32961 (n_15835, n17384);
  and g32962 (n17385, n_15832, n_15835);
  and g32963 (n17386, n_15833, n_15835);
  and g32964 (n17387, n_15834, n17386);
  not g32965 (n_15836, n17385);
  not g32966 (n_15837, n17387);
  and g32967 (n17388, n_15836, n_15837);
  and g32968 (n17389, n17283, n17388);
  not g32969 (n_15838, n17283);
  not g32970 (n_15839, n17388);
  and g32971 (n17390, n_15838, n_15839);
  not g32972 (n_15840, n17389);
  not g32973 (n_15841, n17390);
  and g32974 (n17391, n_15840, n_15841);
  not g32975 (n_15842, n17391);
  and g32976 (n17392, n17281, n_15842);
  not g32977 (n_15843, n17281);
  and g32978 (n17393, n_15843, n_15840);
  and g32979 (n17394, n_15841, n17393);
  not g32980 (n_15844, n17392);
  not g32981 (n_15845, n17394);
  and g32982 (\asquared[103] , n_15844, n_15845);
  not g32983 (n_15846, n17393);
  and g32984 (n17396, n_15841, n_15846);
  and g32985 (n17397, n_15827, n_15834);
  and g32986 (n17398, \a[46] , \a[57] );
  and g32987 (n17399, \a[47] , \a[56] );
  not g32988 (n_15847, n17398);
  not g32989 (n_15848, n17399);
  and g32990 (n17400, n_15847, n_15848);
  and g32991 (n17401, n5666, n8200);
  not g32992 (n_15849, n17401);
  not g32995 (n_15850, n17400);
  not g32997 (n_15851, n17404);
  and g32998 (n17405, n_15849, n_15851);
  and g32999 (n17406, n_15850, n17405);
  and g33000 (n17407, \a[60] , n_15851);
  and g33001 (n17408, \a[43] , n17407);
  not g33002 (n_15852, n17406);
  not g33003 (n_15853, n17408);
  and g33004 (n17409, n_15852, n_15853);
  and g33005 (n17410, n6325, n7699);
  and g33006 (n17411, n5888, n7697);
  and g33007 (n17412, n6256, n7701);
  not g33008 (n_15854, n17411);
  not g33009 (n_15855, n17412);
  and g33010 (n17413, n_15854, n_15855);
  not g33011 (n_15856, n17410);
  not g33012 (n_15857, n17413);
  and g33013 (n17414, n_15856, n_15857);
  not g33014 (n_15858, n17414);
  and g33015 (n17415, \a[55] , n_15858);
  and g33016 (n17416, \a[48] , n17415);
  and g33017 (n17417, n_15856, n_15858);
  and g33018 (n17418, \a[50] , \a[53] );
  not g33019 (n_15859, n12113);
  not g33020 (n_15860, n17418);
  and g33021 (n17419, n_15859, n_15860);
  not g33022 (n_15861, n17419);
  and g33023 (n17420, n17417, n_15861);
  not g33024 (n_15862, n17416);
  not g33025 (n_15863, n17420);
  and g33026 (n17421, n_15862, n_15863);
  not g33027 (n_15864, n17409);
  not g33028 (n_15865, n17421);
  and g33029 (n17422, n_15864, n_15865);
  not g33030 (n_15866, n17422);
  and g33031 (n17423, n_15864, n_15866);
  and g33032 (n17424, n_15865, n_15866);
  not g33033 (n_15867, n17423);
  not g33034 (n_15868, n17424);
  and g33035 (n17425, n_15867, n_15868);
  and g33036 (n17426, \a[52] , n13860);
  not g33037 (n_15869, n17426);
  and g33038 (n17427, n6968, n_15869);
  not g33039 (n_15870, n17427);
  and g33040 (n17428, n6968, n_15870);
  and g33041 (n17429, n_15869, n_15870);
  not g33042 (n_15871, \a[52] );
  not g33043 (n_15872, n13860);
  and g33044 (n17430, n_15871, n_15872);
  not g33045 (n_15873, n17430);
  and g33046 (n17431, n17429, n_15873);
  not g33047 (n_15874, n17428);
  not g33048 (n_15875, n17431);
  and g33049 (n17432, n_15874, n_15875);
  not g33050 (n_15876, n17425);
  not g33051 (n_15877, n17432);
  and g33052 (n17433, n_15876, n_15877);
  not g33053 (n_15878, n17433);
  and g33054 (n17434, n_15876, n_15878);
  and g33055 (n17435, n_15877, n_15878);
  not g33056 (n_15879, n17434);
  not g33057 (n_15880, n17435);
  and g33058 (n17436, n_15879, n_15880);
  and g33059 (n17437, \a[40] , \a[63] );
  not g33060 (n_15881, n17344);
  and g33061 (n17438, n_15881, n17437);
  not g33062 (n_15882, n17437);
  and g33063 (n17439, n17344, n_15882);
  not g33064 (n_15883, n17438);
  not g33065 (n_15884, n17439);
  and g33066 (n17440, n_15883, n_15884);
  not g33067 (n_15885, n17440);
  and g33068 (n17441, n17330, n_15885);
  not g33069 (n_15886, n17330);
  and g33070 (n17442, n_15886, n17440);
  not g33071 (n_15887, n17441);
  not g33072 (n_15888, n17442);
  and g33073 (n17443, n_15887, n_15888);
  and g33074 (n17444, n17296, n17316);
  not g33075 (n_15889, n17296);
  not g33076 (n_15890, n17316);
  and g33077 (n17445, n_15889, n_15890);
  not g33078 (n_15891, n17444);
  not g33079 (n_15892, n17445);
  and g33080 (n17446, n_15891, n_15892);
  and g33081 (n17447, n5713, n8987);
  and g33082 (n17448, n4639, n8905);
  and g33083 (n17449, \a[45] , \a[61] );
  and g33084 (n17450, n17125, n17449);
  not g33085 (n_15893, n17448);
  not g33086 (n_15894, n17450);
  and g33087 (n17451, n_15893, n_15894);
  not g33088 (n_15895, n17447);
  not g33089 (n_15896, n17451);
  and g33090 (n17452, n_15895, n_15896);
  not g33091 (n_15897, n17452);
  and g33092 (n17453, \a[61] , n_15897);
  and g33093 (n17454, \a[42] , n17453);
  and g33094 (n17455, \a[45] , \a[58] );
  not g33095 (n_15898, n16983);
  not g33096 (n_15899, n17455);
  and g33097 (n17456, n_15898, n_15899);
  and g33098 (n17457, n_15895, n_15897);
  not g33099 (n_15900, n17456);
  and g33100 (n17458, n_15900, n17457);
  not g33101 (n_15901, n17454);
  not g33102 (n_15902, n17458);
  and g33103 (n17459, n_15901, n_15902);
  not g33104 (n_15903, n17459);
  and g33105 (n17460, n17446, n_15903);
  not g33106 (n_15904, n17460);
  and g33107 (n17461, n17446, n_15904);
  and g33108 (n17462, n_15903, n_15904);
  not g33109 (n_15905, n17461);
  not g33110 (n_15906, n17462);
  and g33111 (n17463, n_15905, n_15906);
  not g33112 (n_15907, n17443);
  and g33113 (n17464, n_15907, n17463);
  not g33114 (n_15908, n17463);
  and g33115 (n17465, n17443, n_15908);
  not g33116 (n_15909, n17464);
  not g33117 (n_15910, n17465);
  and g33118 (n17466, n_15909, n_15910);
  not g33119 (n_15911, n17436);
  and g33120 (n17467, n_15911, n17466);
  not g33121 (n_15912, n17467);
  and g33122 (n17468, n_15911, n_15912);
  and g33123 (n17469, n17466, n_15912);
  not g33124 (n_15913, n17468);
  not g33125 (n_15914, n17469);
  and g33126 (n17470, n_15913, n_15914);
  not g33127 (n_15915, n17397);
  not g33128 (n_15916, n17470);
  and g33129 (n17471, n_15915, n_15916);
  not g33130 (n_15917, n17471);
  and g33131 (n17472, n_15915, n_15917);
  and g33132 (n17473, n_15916, n_15917);
  not g33133 (n_15918, n17472);
  not g33134 (n_15919, n17473);
  and g33135 (n17474, n_15918, n_15919);
  and g33136 (n17475, n_15745, n_15757);
  and g33137 (n17476, n_15812, n_15816);
  and g33138 (n17477, n17475, n17476);
  not g33139 (n_15920, n17475);
  not g33140 (n_15921, n17476);
  and g33141 (n17478, n_15920, n_15921);
  not g33142 (n_15922, n17477);
  not g33143 (n_15923, n17478);
  and g33144 (n17479, n_15922, n_15923);
  and g33145 (n17480, n_15783, n_15798);
  not g33146 (n_15924, n17479);
  and g33147 (n17481, n_15924, n17480);
  not g33148 (n_15925, n17480);
  and g33149 (n17482, n17479, n_15925);
  not g33150 (n_15926, n17481);
  not g33151 (n_15927, n17482);
  and g33152 (n17483, n_15926, n_15927);
  and g33153 (n17484, n_15763, n_15805);
  and g33154 (n17485, n_15820, n_15824);
  and g33155 (n17486, n17484, n17485);
  not g33156 (n_15928, n17484);
  not g33157 (n_15929, n17485);
  and g33158 (n17487, n_15928, n_15929);
  not g33159 (n_15930, n17486);
  not g33160 (n_15931, n17487);
  and g33161 (n17488, n_15930, n_15931);
  and g33162 (n17489, n17483, n17488);
  not g33163 (n_15932, n17483);
  not g33164 (n_15933, n17488);
  and g33165 (n17490, n_15932, n_15933);
  not g33166 (n_15934, n17489);
  not g33167 (n_15935, n17490);
  and g33168 (n17491, n_15934, n_15935);
  not g33169 (n_15936, n17474);
  and g33170 (n17492, n_15936, n17491);
  not g33171 (n_15937, n17492);
  and g33172 (n17493, n_15936, n_15937);
  and g33173 (n17494, n17491, n_15937);
  not g33174 (n_15938, n17493);
  not g33175 (n_15939, n17494);
  and g33176 (n17495, n_15938, n_15939);
  and g33177 (n17496, n_15806, n_15835);
  not g33178 (n_15940, n17495);
  not g33179 (n_15941, n17496);
  and g33180 (n17497, n_15940, n_15941);
  and g33181 (n17498, n17495, n17496);
  not g33182 (n_15942, n17497);
  not g33183 (n_15943, n17498);
  and g33184 (n17499, n_15942, n_15943);
  not g33185 (n_15944, n17396);
  not g33186 (n_15945, n17499);
  and g33187 (n17500, n_15944, n_15945);
  and g33188 (n17501, n17396, n17499);
  or g33189 (\asquared[104] , n17500, n17501);
  and g33190 (n17503, n_15944, n_15943);
  not g33191 (n_15946, n17503);
  and g33192 (n17504, n_15942, n_15946);
  and g33193 (n17505, n_15917, n_15937);
  and g33194 (n17506, n_15931, n_15934);
  and g33195 (n17507, n17405, n17417);
  not g33196 (n_15947, n17405);
  not g33197 (n_15948, n17417);
  and g33198 (n17508, n_15947, n_15948);
  not g33199 (n_15949, n17507);
  not g33200 (n_15950, n17508);
  and g33201 (n17509, n_15949, n_15950);
  not g33202 (n_15951, n17509);
  and g33203 (n17510, n17457, n_15951);
  not g33204 (n_15952, n17457);
  and g33205 (n17511, n_15952, n17509);
  not g33206 (n_15953, n17510);
  not g33207 (n_15954, n17511);
  and g33208 (n17512, n_15953, n_15954);
  and g33209 (n17513, n_15866, n_15878);
  not g33210 (n_15955, n17512);
  and g33211 (n17514, n_15955, n17513);
  not g33212 (n_15956, n17513);
  and g33213 (n17515, n17512, n_15956);
  not g33214 (n_15957, n17514);
  not g33215 (n_15958, n17515);
  and g33216 (n17516, n_15957, n_15958);
  and g33217 (n17517, \a[43] , \a[61] );
  and g33218 (n17518, \a[45] , \a[59] );
  not g33219 (n_15959, n17517);
  not g33220 (n_15960, n17518);
  and g33221 (n17519, n_15959, n_15960);
  and g33222 (n17520, n4811, n8905);
  and g33223 (n17521, n5296, n9512);
  and g33224 (n17522, n5713, n9509);
  not g33225 (n_15961, n17521);
  not g33226 (n_15962, n17522);
  and g33227 (n17523, n_15961, n_15962);
  not g33228 (n_15963, n17520);
  not g33229 (n_15964, n17523);
  and g33230 (n17524, n_15963, n_15964);
  not g33231 (n_15965, n17524);
  and g33232 (n17525, n_15963, n_15965);
  not g33233 (n_15966, n17519);
  and g33234 (n17526, n_15966, n17525);
  and g33235 (n17527, \a[60] , n_15965);
  and g33236 (n17528, \a[44] , n17527);
  not g33237 (n_15967, n17526);
  not g33238 (n_15968, n17528);
  and g33239 (n17529, n_15967, n_15968);
  and g33240 (n17530, n6252, n8200);
  and g33241 (n17531, n5666, n8436);
  and g33242 (n17532, \a[48] , \a[58] );
  and g33243 (n17533, n17327, n17532);
  not g33244 (n_15969, n17531);
  not g33245 (n_15970, n17533);
  and g33246 (n17534, n_15969, n_15970);
  not g33247 (n_15971, n17530);
  not g33248 (n_15972, n17534);
  and g33249 (n17535, n_15971, n_15972);
  not g33250 (n_15973, n17535);
  and g33251 (n17536, \a[58] , n_15973);
  and g33252 (n17537, \a[46] , n17536);
  and g33253 (n17538, n_15971, n_15973);
  and g33254 (n17539, \a[47] , \a[57] );
  not g33255 (n_15974, n9666);
  not g33256 (n_15975, n17539);
  and g33257 (n17540, n_15974, n_15975);
  not g33258 (n_15976, n17540);
  and g33259 (n17541, n17538, n_15976);
  not g33260 (n_15977, n17537);
  not g33261 (n_15978, n17541);
  and g33262 (n17542, n_15977, n_15978);
  not g33263 (n_15979, n17529);
  not g33264 (n_15980, n17542);
  and g33265 (n17543, n_15979, n_15980);
  not g33266 (n_15981, n17543);
  and g33267 (n17544, n_15979, n_15981);
  and g33268 (n17545, n_15980, n_15981);
  not g33269 (n_15982, n17544);
  not g33270 (n_15983, n17545);
  and g33271 (n17546, n_15982, n_15983);
  and g33272 (n17547, n6564, n7699);
  and g33273 (n17548, n7232, n9801);
  and g33274 (n17549, n6325, n7701);
  not g33275 (n_15984, n17548);
  not g33276 (n_15985, n17549);
  and g33277 (n17550, n_15984, n_15985);
  not g33278 (n_15986, n17547);
  not g33279 (n_15987, n17550);
  and g33280 (n17551, n_15986, n_15987);
  not g33281 (n_15988, n17551);
  and g33282 (n17552, n9801, n_15988);
  and g33283 (n17553, n_15986, n_15988);
  and g33284 (n17554, \a[50] , \a[54] );
  not g33285 (n_15989, n7232);
  not g33286 (n_15990, n17554);
  and g33287 (n17555, n_15989, n_15990);
  not g33288 (n_15991, n17555);
  and g33289 (n17556, n17553, n_15991);
  not g33290 (n_15992, n17552);
  not g33291 (n_15993, n17556);
  and g33292 (n17557, n_15992, n_15993);
  not g33293 (n_15994, n17546);
  not g33294 (n_15995, n17557);
  and g33295 (n17558, n_15994, n_15995);
  not g33296 (n_15996, n17558);
  and g33297 (n17559, n_15994, n_15996);
  and g33298 (n17560, n_15995, n_15996);
  not g33299 (n_15997, n17559);
  not g33300 (n_15998, n17560);
  and g33301 (n17561, n_15997, n_15998);
  not g33302 (n_15999, n17561);
  and g33303 (n17562, n17516, n_15999);
  not g33304 (n_16000, n17516);
  and g33305 (n17563, n_16000, n17561);
  not g33306 (n_16001, n17506);
  not g33307 (n_16002, n17563);
  and g33308 (n17564, n_16001, n_16002);
  not g33309 (n_16003, n17562);
  and g33310 (n17565, n_16003, n17564);
  not g33311 (n_16004, n17565);
  and g33312 (n17566, n_16001, n_16004);
  and g33313 (n17567, n_16002, n_16004);
  and g33314 (n17568, n_16003, n17567);
  not g33315 (n_16005, n17566);
  not g33316 (n_16006, n17568);
  and g33317 (n17569, n_16005, n_16006);
  and g33318 (n17570, n_15910, n_15912);
  and g33319 (n17571, n_15923, n_15927);
  and g33320 (n17572, n17570, n17571);
  not g33321 (n_16007, n17570);
  not g33322 (n_16008, n17571);
  and g33323 (n17573, n_16007, n_16008);
  not g33324 (n_16009, n17572);
  not g33325 (n_16010, n17573);
  and g33326 (n17574, n_16009, n_16010);
  and g33327 (n17575, n_15883, n_15888);
  and g33328 (n17576, n5344, n9792);
  and g33329 (n17577, \a[41] , \a[63] );
  not g33330 (n_16011, n14368);
  not g33331 (n_16012, n17577);
  and g33332 (n17578, n_16011, n_16012);
  not g33333 (n_16013, n17576);
  not g33334 (n_16014, n17578);
  and g33335 (n17579, n_16013, n_16014);
  not g33336 (n_16015, n17429);
  and g33337 (n17580, n_16015, n17579);
  not g33338 (n_16016, n17579);
  and g33339 (n17581, n17429, n_16016);
  not g33340 (n_16017, n17580);
  not g33341 (n_16018, n17581);
  and g33342 (n17582, n_16017, n_16018);
  not g33343 (n_16019, n17582);
  and g33344 (n17583, n17575, n_16019);
  not g33345 (n_16020, n17575);
  and g33346 (n17584, n_16020, n17582);
  not g33347 (n_16021, n17583);
  not g33348 (n_16022, n17584);
  and g33349 (n17585, n_16021, n_16022);
  and g33350 (n17586, n_15892, n_15904);
  not g33351 (n_16023, n17585);
  and g33352 (n17587, n_16023, n17586);
  not g33353 (n_16024, n17586);
  and g33354 (n17588, n17585, n_16024);
  not g33355 (n_16025, n17587);
  not g33356 (n_16026, n17588);
  and g33357 (n17589, n_16025, n_16026);
  and g33358 (n17590, n17574, n17589);
  not g33359 (n_16027, n17574);
  not g33360 (n_16028, n17589);
  and g33361 (n17591, n_16027, n_16028);
  not g33362 (n_16029, n17590);
  not g33363 (n_16030, n17591);
  and g33364 (n17592, n_16029, n_16030);
  not g33365 (n_16031, n17569);
  and g33366 (n17593, n_16031, n17592);
  not g33367 (n_16032, n17593);
  and g33368 (n17594, n_16031, n_16032);
  and g33369 (n17595, n17592, n_16032);
  not g33370 (n_16033, n17594);
  not g33371 (n_16034, n17595);
  and g33372 (n17596, n_16033, n_16034);
  not g33373 (n_16035, n17505);
  not g33374 (n_16036, n17596);
  and g33375 (n17597, n_16035, n_16036);
  and g33376 (n17598, n17505, n17596);
  not g33377 (n_16037, n17597);
  not g33378 (n_16038, n17598);
  and g33379 (n17599, n_16037, n_16038);
  not g33380 (n_16039, n17504);
  and g33381 (n17600, n_16039, n17599);
  not g33382 (n_16040, n17599);
  and g33383 (n17601, n17504, n_16040);
  not g33384 (n_16041, n17600);
  not g33385 (n_16042, n17601);
  and g33386 (\asquared[105] , n_16041, n_16042);
  and g33387 (n17603, n17538, n17553);
  not g33388 (n_16043, n17538);
  not g33389 (n_16044, n17553);
  and g33390 (n17604, n_16043, n_16044);
  not g33391 (n_16045, n17603);
  not g33392 (n_16046, n17604);
  and g33393 (n17605, n_16045, n_16046);
  not g33394 (n_16047, n17605);
  and g33395 (n17606, n17525, n_16047);
  not g33396 (n_16048, n17525);
  and g33397 (n17607, n_16048, n17605);
  not g33398 (n_16049, n17606);
  not g33399 (n_16050, n17607);
  and g33400 (n17608, n_16049, n_16050);
  and g33401 (n17609, n_15981, n_15996);
  not g33402 (n_16051, n17608);
  and g33403 (n17610, n_16051, n17609);
  not g33404 (n_16052, n17609);
  and g33405 (n17611, n17608, n_16052);
  not g33406 (n_16053, n17610);
  not g33407 (n_16054, n17611);
  and g33408 (n17612, n_16053, n_16054);
  and g33409 (n17613, n_16022, n_16026);
  not g33410 (n_16055, n17612);
  and g33411 (n17614, n_16055, n17613);
  not g33412 (n_16056, n17613);
  and g33413 (n17615, n17612, n_16056);
  not g33414 (n_16057, n17614);
  not g33415 (n_16058, n17615);
  and g33416 (n17616, n_16057, n_16058);
  and g33417 (n17617, n_16010, n_16029);
  not g33418 (n_16059, n17617);
  and g33419 (n17618, n17616, n_16059);
  not g33420 (n_16060, n17616);
  and g33421 (n17619, n_16060, n17617);
  not g33422 (n_16061, n17618);
  not g33423 (n_16062, n17619);
  and g33424 (n17620, n_16061, n_16062);
  and g33425 (n17621, n_15958, n_16003);
  and g33426 (n17622, \a[62] , n16612);
  not g33427 (n_16063, n17622);
  and g33428 (n17623, n7433, n_16063);
  not g33429 (n_16064, n17623);
  and g33430 (n17624, n_16063, n_16064);
  not g33431 (n_16065, \a[53] );
  not g33432 (n_16066, n14732);
  and g33433 (n17625, n_16065, n_16066);
  not g33434 (n_16067, n17625);
  and g33435 (n17626, n17624, n_16067);
  and g33436 (n17627, n7433, n_16064);
  not g33437 (n_16068, n17626);
  not g33438 (n_16069, n17627);
  and g33439 (n17628, n_16068, n_16069);
  and g33440 (n17629, n6564, n7701);
  and g33441 (n17630, n7421, n9934);
  and g33442 (n17631, n6325, n9161);
  not g33443 (n_16070, n17630);
  not g33444 (n_16071, n17631);
  and g33445 (n17632, n_16070, n_16071);
  not g33446 (n_16072, n17629);
  not g33447 (n_16073, n17632);
  and g33448 (n17633, n_16072, n_16073);
  not g33449 (n_16074, n17633);
  and g33450 (n17634, \a[56] , n_16074);
  and g33451 (n17635, \a[49] , n17634);
  and g33452 (n17636, \a[51] , \a[54] );
  and g33453 (n17637, \a[50] , \a[55] );
  not g33454 (n_16075, n17636);
  not g33455 (n_16076, n17637);
  and g33456 (n17638, n_16075, n_16076);
  and g33457 (n17639, n_16072, n_16074);
  not g33458 (n_16077, n17638);
  and g33459 (n17640, n_16077, n17639);
  not g33460 (n_16078, n17635);
  not g33461 (n_16079, n17640);
  and g33462 (n17641, n_16078, n_16079);
  not g33463 (n_16080, n17628);
  not g33464 (n_16081, n17641);
  and g33465 (n17642, n_16080, n_16081);
  not g33466 (n_16082, n17642);
  and g33467 (n17643, n_16080, n_16082);
  and g33468 (n17644, n_16081, n_16082);
  not g33469 (n_16083, n17643);
  not g33470 (n_16084, n17644);
  and g33471 (n17645, n_16083, n_16084);
  and g33472 (n17646, n_15950, n_15954);
  and g33473 (n17647, n17645, n17646);
  not g33474 (n_16085, n17645);
  not g33475 (n_16086, n17646);
  and g33476 (n17648, n_16085, n_16086);
  not g33477 (n_16087, n17647);
  not g33478 (n_16088, n17648);
  and g33479 (n17649, n_16087, n_16088);
  and g33480 (n17650, n5713, n9512);
  and g33481 (n17651, n11634, n15167);
  and g33482 (n17652, n4639, n9909);
  not g33483 (n_16089, n17651);
  not g33484 (n_16090, n17652);
  and g33485 (n17653, n_16089, n_16090);
  not g33486 (n_16091, n17650);
  not g33487 (n_16092, n17653);
  and g33488 (n17654, n_16091, n_16092);
  not g33489 (n_16093, n17654);
  and g33490 (n17655, \a[42] , n_16093);
  and g33491 (n17656, \a[63] , n17655);
  and g33492 (n17657, n_16091, n_16093);
  and g33493 (n17658, \a[44] , \a[61] );
  and g33494 (n17659, \a[45] , \a[60] );
  not g33495 (n_16094, n17658);
  not g33496 (n_16095, n17659);
  and g33497 (n17660, n_16094, n_16095);
  not g33498 (n_16096, n17660);
  and g33499 (n17661, n17657, n_16096);
  not g33500 (n_16097, n17656);
  not g33501 (n_16098, n17661);
  and g33502 (n17662, n_16097, n_16098);
  and g33503 (n17663, n_16013, n_16017);
  not g33504 (n_16099, n17662);
  and g33505 (n17664, n_16099, n17663);
  not g33506 (n_16100, n17663);
  and g33507 (n17665, n17662, n_16100);
  not g33508 (n_16101, n17664);
  not g33509 (n_16102, n17665);
  and g33510 (n17666, n_16101, n_16102);
  and g33511 (n17667, n6252, n8436);
  and g33512 (n17668, n8578, n8985);
  and g33513 (n17669, n5666, n8987);
  not g33514 (n_16103, n17668);
  not g33515 (n_16104, n17669);
  and g33516 (n17670, n_16103, n_16104);
  not g33517 (n_16105, n17667);
  not g33518 (n_16106, n17670);
  and g33519 (n17671, n_16105, n_16106);
  not g33520 (n_16107, n17671);
  and g33521 (n17672, \a[59] , n_16107);
  and g33522 (n17673, \a[46] , n17672);
  and g33523 (n17674, n_16105, n_16107);
  and g33524 (n17675, \a[47] , \a[58] );
  and g33525 (n17676, \a[48] , \a[57] );
  not g33526 (n_16108, n17675);
  not g33527 (n_16109, n17676);
  and g33528 (n17677, n_16108, n_16109);
  not g33529 (n_16110, n17677);
  and g33530 (n17678, n17674, n_16110);
  not g33531 (n_16111, n17673);
  not g33532 (n_16112, n17678);
  and g33533 (n17679, n_16111, n_16112);
  not g33534 (n_16113, n17666);
  not g33535 (n_16114, n17679);
  and g33536 (n17680, n_16113, n_16114);
  and g33537 (n17681, n17666, n17679);
  not g33538 (n_16115, n17680);
  not g33539 (n_16116, n17681);
  and g33540 (n17682, n_16115, n_16116);
  not g33541 (n_16117, n17649);
  not g33542 (n_16118, n17682);
  and g33543 (n17683, n_16117, n_16118);
  and g33544 (n17684, n17649, n17682);
  not g33545 (n_16119, n17683);
  not g33546 (n_16120, n17684);
  and g33547 (n17685, n_16119, n_16120);
  not g33548 (n_16121, n17621);
  and g33549 (n17686, n_16121, n17685);
  not g33550 (n_16122, n17685);
  and g33551 (n17687, n17621, n_16122);
  not g33552 (n_16123, n17686);
  not g33553 (n_16124, n17687);
  and g33554 (n17688, n_16123, n_16124);
  and g33555 (n17689, n17620, n17688);
  not g33556 (n_16125, n17620);
  not g33557 (n_16126, n17688);
  and g33558 (n17690, n_16125, n_16126);
  not g33559 (n_16127, n17689);
  not g33560 (n_16128, n17690);
  and g33561 (n17691, n_16127, n_16128);
  and g33562 (n17692, n_16004, n_16032);
  not g33563 (n_16129, n17691);
  and g33564 (n17693, n_16129, n17692);
  not g33565 (n_16130, n17692);
  and g33566 (n17694, n17691, n_16130);
  not g33567 (n_16131, n17693);
  not g33568 (n_16132, n17694);
  and g33569 (n17695, n_16131, n_16132);
  and g33570 (n17696, n_16039, n_16038);
  not g33571 (n_16133, n17696);
  and g33572 (n17697, n_16037, n_16133);
  not g33573 (n_16134, n17695);
  and g33574 (n17698, n_16134, n17697);
  not g33575 (n_16135, n17697);
  and g33576 (n17699, n17695, n_16135);
  not g33577 (n_16136, n17698);
  not g33578 (n_16137, n17699);
  and g33579 (\asquared[106] , n_16136, n_16137);
  and g33580 (n17701, n_16131, n_16135);
  not g33581 (n_16138, n17701);
  and g33582 (n17702, n_16132, n_16138);
  and g33583 (n17703, n_16061, n_16127);
  and g33584 (n17704, n_16054, n_16058);
  and g33585 (n17705, n6256, n8436);
  and g33586 (n17706, n6254, n8985);
  and g33587 (n17707, n6252, n8987);
  not g33588 (n_16139, n17706);
  not g33589 (n_16140, n17707);
  and g33590 (n17708, n_16139, n_16140);
  not g33591 (n_16141, n17705);
  not g33592 (n_16142, n17708);
  and g33593 (n17709, n_16141, n_16142);
  not g33594 (n_16143, n17709);
  and g33595 (n17710, n_16141, n_16143);
  not g33596 (n_16144, n12601);
  not g33597 (n_16145, n17532);
  and g33598 (n17711, n_16144, n_16145);
  not g33599 (n_16146, n17711);
  and g33600 (n17712, n17710, n_16146);
  and g33601 (n17713, \a[59] , n_16143);
  and g33602 (n17714, \a[47] , n17713);
  not g33603 (n_16147, n17712);
  not g33604 (n_16148, n17714);
  and g33605 (n17715, n_16147, n_16148);
  and g33606 (n17716, n6968, n7701);
  and g33607 (n17717, n6966, n7421);
  and g33608 (n17718, n6564, n9161);
  not g33609 (n_16149, n17717);
  not g33610 (n_16150, n17718);
  and g33611 (n17719, n_16149, n_16150);
  not g33612 (n_16151, n17716);
  not g33613 (n_16152, n17719);
  and g33614 (n17720, n_16151, n_16152);
  not g33615 (n_16153, n17720);
  and g33616 (n17721, \a[56] , n_16153);
  and g33617 (n17722, \a[50] , n17721);
  and g33618 (n17723, n_16151, n_16153);
  and g33619 (n17724, \a[51] , \a[55] );
  not g33620 (n_16154, n10905);
  not g33621 (n_16155, n17724);
  and g33622 (n17725, n_16154, n_16155);
  not g33623 (n_16156, n17725);
  and g33624 (n17726, n17723, n_16156);
  not g33625 (n_16157, n17722);
  not g33626 (n_16158, n17726);
  and g33627 (n17727, n_16157, n_16158);
  not g33628 (n_16159, n17715);
  not g33629 (n_16160, n17727);
  and g33630 (n17728, n_16159, n_16160);
  not g33631 (n_16161, n17728);
  and g33632 (n17729, n_16159, n_16161);
  and g33633 (n17730, n_16160, n_16161);
  not g33634 (n_16162, n17729);
  not g33635 (n_16163, n17730);
  and g33636 (n17731, n_16162, n_16163);
  and g33637 (n17732, n_16046, n_16050);
  and g33638 (n17733, n17731, n17732);
  not g33639 (n_16164, n17731);
  not g33640 (n_16165, n17732);
  and g33641 (n17734, n_16164, n_16165);
  not g33642 (n_16166, n17733);
  not g33643 (n_16167, n17734);
  and g33644 (n17735, n_16166, n_16167);
  and g33645 (n17736, n17657, n17674);
  not g33646 (n_16168, n17657);
  not g33647 (n_16169, n17674);
  and g33648 (n17737, n_16168, n_16169);
  not g33649 (n_16170, n17736);
  not g33650 (n_16171, n17737);
  and g33651 (n17738, n_16170, n_16171);
  and g33652 (n17739, n5560, n9512);
  and g33653 (n17740, n5713, n9721);
  and g33654 (n17741, \a[46] , \a[60] );
  and g33655 (n17742, n15107, n17741);
  not g33656 (n_16172, n17740);
  not g33657 (n_16173, n17742);
  and g33658 (n17743, n_16172, n_16173);
  not g33659 (n_16174, n17739);
  not g33660 (n_16175, n17743);
  and g33661 (n17744, n_16174, n_16175);
  not g33662 (n_16176, n17744);
  and g33663 (n17745, n15107, n_16176);
  and g33664 (n17746, n_16174, n_16176);
  not g33665 (n_16177, n17449);
  not g33666 (n_16178, n17741);
  and g33667 (n17747, n_16177, n_16178);
  not g33668 (n_16179, n17747);
  and g33669 (n17748, n17746, n_16179);
  not g33670 (n_16180, n17745);
  not g33671 (n_16181, n17748);
  and g33672 (n17749, n_16180, n_16181);
  not g33673 (n_16182, n17749);
  and g33674 (n17750, n17738, n_16182);
  not g33675 (n_16183, n17750);
  and g33676 (n17751, n17738, n_16183);
  and g33677 (n17752, n_16182, n_16183);
  not g33678 (n_16184, n17751);
  not g33679 (n_16185, n17752);
  and g33680 (n17753, n_16184, n_16185);
  not g33681 (n_16186, n17753);
  and g33682 (n17754, n17735, n_16186);
  not g33683 (n_16187, n17735);
  and g33684 (n17755, n_16187, n17753);
  not g33685 (n_16188, n17704);
  not g33686 (n_16189, n17755);
  and g33687 (n17756, n_16188, n_16189);
  not g33688 (n_16190, n17754);
  and g33689 (n17757, n_16190, n17756);
  not g33690 (n_16191, n17757);
  and g33691 (n17758, n_16188, n_16191);
  and g33692 (n17759, n_16190, n_16191);
  and g33693 (n17760, n_16189, n17759);
  not g33694 (n_16192, n17758);
  not g33695 (n_16193, n17760);
  and g33696 (n17761, n_16192, n_16193);
  and g33697 (n17762, \a[43] , \a[63] );
  not g33698 (n_16194, n17624);
  and g33699 (n17763, n_16194, n17762);
  not g33700 (n_16195, n17762);
  and g33701 (n17764, n17624, n_16195);
  not g33702 (n_16196, n17763);
  not g33703 (n_16197, n17764);
  and g33704 (n17765, n_16196, n_16197);
  not g33705 (n_16198, n17765);
  and g33706 (n17766, n17639, n_16198);
  not g33707 (n_16199, n17639);
  and g33708 (n17767, n_16199, n17765);
  not g33709 (n_16200, n17766);
  not g33710 (n_16201, n17767);
  and g33711 (n17768, n_16200, n_16201);
  and g33712 (n17769, n_16099, n_16100);
  not g33713 (n_16202, n17769);
  and g33714 (n17770, n_16115, n_16202);
  not g33715 (n_16203, n17768);
  and g33716 (n17771, n_16203, n17770);
  not g33717 (n_16204, n17770);
  and g33718 (n17772, n17768, n_16204);
  not g33719 (n_16205, n17771);
  not g33720 (n_16206, n17772);
  and g33721 (n17773, n_16205, n_16206);
  and g33722 (n17774, n_16082, n_16088);
  not g33723 (n_16207, n17773);
  and g33724 (n17775, n_16207, n17774);
  not g33725 (n_16208, n17774);
  and g33726 (n17776, n17773, n_16208);
  not g33727 (n_16209, n17775);
  not g33728 (n_16210, n17776);
  and g33729 (n17777, n_16209, n_16210);
  and g33730 (n17778, n_16120, n_16123);
  not g33731 (n_16211, n17778);
  and g33732 (n17779, n17777, n_16211);
  not g33733 (n_16212, n17777);
  and g33734 (n17780, n_16212, n17778);
  not g33735 (n_16213, n17779);
  not g33736 (n_16214, n17780);
  and g33737 (n17781, n_16213, n_16214);
  and g33738 (n17782, n17761, n17781);
  not g33739 (n_16215, n17761);
  not g33740 (n_16216, n17781);
  and g33741 (n17783, n_16215, n_16216);
  not g33742 (n_16217, n17782);
  not g33743 (n_16218, n17783);
  and g33744 (n17784, n_16217, n_16218);
  not g33745 (n_16219, n17703);
  not g33746 (n_16220, n17784);
  and g33747 (n17785, n_16219, n_16220);
  and g33748 (n17786, n17703, n17784);
  not g33749 (n_16221, n17785);
  not g33750 (n_16222, n17786);
  and g33751 (n17787, n_16221, n_16222);
  not g33752 (n_16223, n17787);
  and g33753 (n17788, n17702, n_16223);
  not g33754 (n_16224, n17702);
  and g33755 (n17789, n_16224, n_16222);
  and g33756 (n17790, n_16221, n17789);
  not g33757 (n_16225, n17788);
  not g33758 (n_16226, n17790);
  and g33759 (\asquared[107] , n_16225, n_16226);
  not g33760 (n_16227, n17789);
  and g33761 (n17792, n_16221, n_16227);
  and g33762 (n17793, n_16215, n17781);
  not g33763 (n_16228, n17793);
  and g33764 (n17794, n_16213, n_16228);
  and g33765 (n17795, n_16206, n_16210);
  and g33766 (n17796, n17710, n17746);
  not g33767 (n_16229, n17710);
  not g33768 (n_16230, n17746);
  and g33769 (n17797, n_16229, n_16230);
  not g33770 (n_16231, n17796);
  not g33771 (n_16232, n17797);
  and g33772 (n17798, n_16231, n_16232);
  and g33773 (n17799, \a[58] , \a[63] );
  and g33774 (n17800, n8252, n17799);
  and g33775 (n17801, n6256, n8987);
  and g33776 (n17802, \a[59] , \a[63] );
  and g33777 (n17803, n15979, n17802);
  not g33778 (n_16233, n17801);
  not g33779 (n_16234, n17803);
  and g33780 (n17804, n_16233, n_16234);
  not g33781 (n_16235, n17800);
  not g33782 (n_16236, n17804);
  and g33783 (n17805, n_16235, n_16236);
  not g33784 (n_16237, n17805);
  and g33785 (n17806, \a[59] , n_16237);
  and g33786 (n17807, \a[48] , n17806);
  and g33787 (n17808, \a[44] , \a[63] );
  and g33788 (n17809, \a[49] , \a[58] );
  not g33789 (n_16238, n17808);
  not g33790 (n_16239, n17809);
  and g33791 (n17810, n_16238, n_16239);
  and g33792 (n17811, n_16235, n_16237);
  not g33793 (n_16240, n17810);
  and g33794 (n17812, n_16240, n17811);
  not g33795 (n_16241, n17807);
  not g33796 (n_16242, n17812);
  and g33797 (n17813, n_16241, n_16242);
  not g33798 (n_16243, n17813);
  and g33799 (n17814, n17798, n_16243);
  not g33800 (n_16244, n17814);
  and g33801 (n17815, n17798, n_16244);
  and g33802 (n17816, n_16243, n_16244);
  not g33803 (n_16245, n17815);
  not g33804 (n_16246, n17816);
  and g33805 (n17817, n_16245, n_16246);
  and g33806 (n17818, \a[54] , n15463);
  not g33807 (n_16247, n17818);
  and g33808 (n17819, n7699, n_16247);
  not g33809 (n_16248, n17819);
  and g33810 (n17820, n_16247, n_16248);
  not g33811 (n_16249, \a[54] );
  not g33812 (n_16250, n15463);
  and g33813 (n17821, n_16249, n_16250);
  not g33814 (n_16251, n17821);
  and g33815 (n17822, n17820, n_16251);
  and g33816 (n17823, n7699, n_16248);
  not g33817 (n_16252, n17822);
  not g33818 (n_16253, n17823);
  and g33819 (n17824, n_16252, n_16253);
  and g33820 (n17825, n6968, n9161);
  and g33821 (n17826, n6966, n11718);
  and g33822 (n17827, n6564, n8200);
  not g33823 (n_16254, n17826);
  not g33824 (n_16255, n17827);
  and g33825 (n17828, n_16254, n_16255);
  not g33826 (n_16256, n17825);
  not g33827 (n_16257, n17828);
  and g33828 (n17829, n_16256, n_16257);
  not g33829 (n_16258, n17829);
  and g33830 (n17830, \a[57] , n_16258);
  and g33831 (n17831, \a[50] , n17830);
  and g33832 (n17832, n_16256, n_16258);
  and g33833 (n17833, \a[51] , \a[56] );
  not g33834 (n_16259, n12388);
  not g33835 (n_16260, n17833);
  and g33836 (n17834, n_16259, n_16260);
  not g33837 (n_16261, n17834);
  and g33838 (n17835, n17832, n_16261);
  not g33839 (n_16262, n17831);
  not g33840 (n_16263, n17835);
  and g33841 (n17836, n_16262, n_16263);
  not g33842 (n_16264, n17824);
  not g33843 (n_16265, n17836);
  and g33844 (n17837, n_16264, n_16265);
  not g33845 (n_16266, n17837);
  and g33846 (n17838, n_16264, n_16266);
  and g33847 (n17839, n_16265, n_16266);
  not g33848 (n_16267, n17838);
  not g33849 (n_16268, n17839);
  and g33850 (n17840, n_16267, n_16268);
  and g33851 (n17841, n5666, n9512);
  not g33852 (n_16269, n17841);
  and g33853 (n17842, \a[60] , n_16269);
  and g33854 (n17843, \a[47] , n17842);
  and g33855 (n17844, \a[46] , n_16269);
  and g33856 (n17845, \a[61] , n17844);
  not g33857 (n_16270, n17843);
  not g33858 (n_16271, n17845);
  and g33859 (n17846, n_16270, n_16271);
  not g33860 (n_16272, n17723);
  not g33861 (n_16273, n17846);
  and g33862 (n17847, n_16272, n_16273);
  not g33863 (n_16274, n17847);
  and g33864 (n17848, n_16272, n_16274);
  and g33865 (n17849, n_16273, n_16274);
  not g33866 (n_16275, n17848);
  not g33867 (n_16276, n17849);
  and g33868 (n17850, n_16275, n_16276);
  not g33869 (n_16277, n17840);
  and g33870 (n17851, n_16277, n17850);
  not g33871 (n_16278, n17850);
  and g33872 (n17852, n17840, n_16278);
  not g33873 (n_16279, n17851);
  not g33874 (n_16280, n17852);
  and g33875 (n17853, n_16279, n_16280);
  not g33876 (n_16281, n17817);
  not g33877 (n_16282, n17853);
  and g33878 (n17854, n_16281, n_16282);
  and g33879 (n17855, n17817, n17853);
  not g33880 (n_16283, n17854);
  not g33881 (n_16284, n17855);
  and g33882 (n17856, n_16283, n_16284);
  not g33883 (n_16285, n17856);
  and g33884 (n17857, n17795, n_16285);
  not g33885 (n_16286, n17795);
  and g33886 (n17858, n_16286, n17856);
  not g33887 (n_16287, n17857);
  not g33888 (n_16288, n17858);
  and g33889 (n17859, n_16287, n_16288);
  and g33890 (n17860, n_16171, n_16183);
  and g33891 (n17861, n_16196, n_16201);
  and g33892 (n17862, n17860, n17861);
  not g33893 (n_16289, n17860);
  not g33894 (n_16290, n17861);
  and g33895 (n17863, n_16289, n_16290);
  not g33896 (n_16291, n17862);
  not g33897 (n_16292, n17863);
  and g33898 (n17864, n_16291, n_16292);
  and g33899 (n17865, n_16161, n_16167);
  not g33900 (n_16293, n17864);
  and g33901 (n17866, n_16293, n17865);
  not g33902 (n_16294, n17865);
  and g33903 (n17867, n17864, n_16294);
  not g33904 (n_16295, n17866);
  not g33905 (n_16296, n17867);
  and g33906 (n17868, n_16295, n_16296);
  not g33907 (n_16297, n17759);
  and g33908 (n17869, n_16297, n17868);
  not g33909 (n_16298, n17868);
  and g33910 (n17870, n17759, n_16298);
  not g33911 (n_16299, n17869);
  not g33912 (n_16300, n17870);
  and g33913 (n17871, n_16299, n_16300);
  and g33914 (n17872, n17859, n17871);
  not g33915 (n_16301, n17859);
  not g33916 (n_16302, n17871);
  and g33917 (n17873, n_16301, n_16302);
  not g33918 (n_16303, n17872);
  not g33919 (n_16304, n17873);
  and g33920 (n17874, n_16303, n_16304);
  not g33921 (n_16305, n17874);
  and g33922 (n17875, n17794, n_16305);
  not g33923 (n_16306, n17794);
  and g33924 (n17876, n_16306, n17874);
  not g33925 (n_16307, n17875);
  not g33926 (n_16308, n17876);
  and g33927 (n17877, n_16307, n_16308);
  not g33928 (n_16309, n17792);
  not g33929 (n_16310, n17877);
  and g33930 (n17878, n_16309, n_16310);
  and g33931 (n17879, n17792, n17877);
  or g33932 (\asquared[108] , n17878, n17879);
  and g33933 (n17881, n_16309, n_16307);
  not g33934 (n_16311, n17881);
  and g33935 (n17882, n_16308, n_16311);
  and g33936 (n17883, n_16299, n_16303);
  and g33937 (n17884, n_16232, n_16244);
  and g33938 (n17885, n7433, n9161);
  and g33939 (n17886, n7232, n11718);
  and g33940 (n17887, n6968, n8200);
  not g33941 (n_16312, n17886);
  not g33942 (n_16313, n17887);
  and g33943 (n17888, n_16312, n_16313);
  not g33944 (n_16314, n17885);
  not g33945 (n_16315, n17888);
  and g33946 (n17889, n_16314, n_16315);
  not g33947 (n_16316, n17889);
  and g33948 (n17890, n14417, n_16316);
  and g33949 (n17891, n_16314, n_16316);
  and g33950 (n17892, \a[52] , \a[56] );
  not g33951 (n_16317, n7697);
  not g33952 (n_16318, n17892);
  and g33953 (n17893, n_16317, n_16318);
  not g33954 (n_16319, n17893);
  and g33955 (n17894, n17891, n_16319);
  not g33956 (n_16320, n17890);
  not g33957 (n_16321, n17894);
  and g33958 (n17895, n_16320, n_16321);
  not g33959 (n_16322, n17884);
  not g33960 (n_16323, n17895);
  and g33961 (n17896, n_16322, n_16323);
  not g33962 (n_16324, n17896);
  and g33963 (n17897, n_16322, n_16324);
  and g33964 (n17898, n_16323, n_16324);
  not g33965 (n_16325, n17897);
  not g33966 (n_16326, n17898);
  and g33967 (n17899, n_16325, n_16326);
  and g33968 (n17900, n_16277, n_16278);
  not g33969 (n_16327, n17900);
  and g33970 (n17901, n_16266, n_16327);
  not g33971 (n_16328, n17899);
  not g33972 (n_16329, n17901);
  and g33973 (n17902, n_16328, n_16329);
  not g33974 (n_16330, n17902);
  and g33975 (n17903, n_16328, n_16330);
  and g33976 (n17904, n_16329, n_16330);
  not g33977 (n_16331, n17903);
  not g33978 (n_16332, n17904);
  and g33979 (n17905, n_16331, n_16332);
  and g33980 (n17906, n_16283, n_16288);
  and g33981 (n17907, n17905, n17906);
  not g33982 (n_16333, n17905);
  not g33983 (n_16334, n17906);
  and g33984 (n17908, n_16333, n_16334);
  not g33985 (n_16335, n17907);
  not g33986 (n_16336, n17908);
  and g33987 (n17909, n_16335, n_16336);
  and g33988 (n17910, n17820, n17832);
  not g33989 (n_16337, n17820);
  not g33990 (n_16338, n17832);
  and g33991 (n17911, n_16337, n_16338);
  not g33992 (n_16339, n17910);
  not g33993 (n_16340, n17911);
  and g33994 (n17912, n_16339, n_16340);
  not g33995 (n_16341, n17912);
  and g33996 (n17913, n17811, n_16341);
  not g33997 (n_16342, n17811);
  and g33998 (n17914, n_16342, n17912);
  not g33999 (n_16343, n17913);
  not g34000 (n_16344, n17914);
  and g34001 (n17915, n_16343, n_16344);
  and g34002 (n17916, n_16292, n_16296);
  not g34003 (n_16345, n17915);
  and g34004 (n17917, n_16345, n17916);
  not g34005 (n_16346, n17916);
  and g34006 (n17918, n17915, n_16346);
  not g34007 (n_16347, n17917);
  not g34008 (n_16348, n17918);
  and g34009 (n17919, n_16347, n_16348);
  and g34010 (n17920, n5666, n9721);
  and g34011 (n17921, n5250, n9909);
  and g34012 (n17922, n5560, n9792);
  not g34013 (n_16349, n17921);
  not g34014 (n_16350, n17922);
  and g34015 (n17923, n_16349, n_16350);
  not g34016 (n_16351, n17920);
  not g34017 (n_16352, n17923);
  and g34018 (n17924, n_16351, n_16352);
  not g34019 (n_16353, n17924);
  and g34020 (n17925, \a[45] , n_16353);
  and g34021 (n17926, \a[63] , n17925);
  and g34022 (n17927, n_16351, n_16353);
  and g34023 (n17928, \a[47] , \a[61] );
  not g34024 (n_16354, n15856);
  not g34025 (n_16355, n17928);
  and g34026 (n17929, n_16354, n_16355);
  not g34027 (n_16356, n17929);
  and g34028 (n17930, n17927, n_16356);
  not g34029 (n_16357, n17926);
  not g34030 (n_16358, n17930);
  and g34031 (n17931, n_16357, n_16358);
  and g34032 (n17932, n_16269, n_16274);
  not g34033 (n_16359, n17931);
  and g34034 (n17933, n_16359, n17932);
  not g34035 (n_16360, n17932);
  and g34036 (n17934, n17931, n_16360);
  not g34037 (n_16361, n17933);
  not g34038 (n_16362, n17934);
  and g34039 (n17935, n_16361, n_16362);
  and g34040 (n17936, n6325, n8987);
  and g34041 (n17937, n5888, n10089);
  and g34042 (n17938, n6256, n9509);
  not g34043 (n_16363, n17937);
  not g34044 (n_16364, n17938);
  and g34045 (n17939, n_16363, n_16364);
  not g34046 (n_16365, n17936);
  not g34047 (n_16366, n17939);
  and g34048 (n17940, n_16365, n_16366);
  not g34049 (n_16367, n17940);
  and g34050 (n17941, \a[60] , n_16367);
  and g34051 (n17942, \a[48] , n17941);
  and g34052 (n17943, \a[49] , \a[59] );
  and g34053 (n17944, \a[50] , \a[58] );
  not g34054 (n_16368, n17943);
  not g34055 (n_16369, n17944);
  and g34056 (n17945, n_16368, n_16369);
  and g34057 (n17946, n_16365, n_16367);
  not g34058 (n_16370, n17945);
  and g34059 (n17947, n_16370, n17946);
  not g34060 (n_16371, n17942);
  not g34061 (n_16372, n17947);
  and g34062 (n17948, n_16371, n_16372);
  not g34063 (n_16373, n17935);
  not g34064 (n_16374, n17948);
  and g34065 (n17949, n_16373, n_16374);
  and g34066 (n17950, n17935, n17948);
  not g34067 (n_16375, n17949);
  not g34068 (n_16376, n17950);
  and g34069 (n17951, n_16375, n_16376);
  and g34070 (n17952, n17919, n17951);
  not g34071 (n_16377, n17919);
  not g34072 (n_16378, n17951);
  and g34073 (n17953, n_16377, n_16378);
  not g34074 (n_16379, n17953);
  and g34075 (n17954, n17909, n_16379);
  not g34076 (n_16380, n17952);
  and g34077 (n17955, n_16380, n17954);
  not g34078 (n_16381, n17955);
  and g34079 (n17956, n17909, n_16381);
  and g34080 (n17957, n_16379, n_16381);
  and g34081 (n17958, n_16380, n17957);
  not g34082 (n_16382, n17956);
  not g34083 (n_16383, n17958);
  and g34084 (n17959, n_16382, n_16383);
  and g34085 (n17960, n17883, n17959);
  not g34086 (n_16384, n17883);
  not g34087 (n_16385, n17959);
  and g34088 (n17961, n_16384, n_16385);
  not g34089 (n_16386, n17960);
  not g34090 (n_16387, n17961);
  and g34091 (n17962, n_16386, n_16387);
  not g34092 (n_16388, n17962);
  and g34093 (n17963, n17882, n_16388);
  not g34094 (n_16389, n17882);
  and g34095 (n17964, n_16389, n_16386);
  and g34096 (n17965, n_16387, n17964);
  not g34097 (n_16390, n17963);
  not g34098 (n_16391, n17965);
  and g34099 (\asquared[109] , n_16390, n_16391);
  not g34100 (n_16392, n17964);
  and g34101 (n17967, n_16387, n_16392);
  and g34102 (n17968, n_16340, n_16344);
  and g34103 (n17969, \a[55] , n16194);
  not g34104 (n_16393, n17969);
  and g34105 (n17970, n7701, n_16393);
  not g34106 (n_16394, n17970);
  and g34107 (n17971, n7701, n_16394);
  and g34108 (n17972, n_16393, n_16394);
  not g34109 (n_16395, \a[55] );
  not g34110 (n_16396, n16194);
  and g34111 (n17973, n_16395, n_16396);
  not g34112 (n_16397, n17973);
  and g34113 (n17974, n17972, n_16397);
  not g34114 (n_16398, n17971);
  not g34115 (n_16399, n17974);
  and g34116 (n17975, n_16398, n_16399);
  not g34117 (n_16400, n17968);
  not g34118 (n_16401, n17975);
  and g34119 (n17976, n_16400, n_16401);
  not g34120 (n_16402, n17976);
  and g34121 (n17977, n_16400, n_16402);
  and g34122 (n17978, n_16401, n_16402);
  not g34123 (n_16403, n17977);
  not g34124 (n_16404, n17978);
  and g34125 (n17979, n_16403, n_16404);
  and g34126 (n17980, n_16359, n_16360);
  not g34127 (n_16405, n17980);
  and g34128 (n17981, n_16375, n_16405);
  and g34129 (n17982, n17979, n17981);
  not g34130 (n_16406, n17979);
  not g34131 (n_16407, n17981);
  and g34132 (n17983, n_16406, n_16407);
  not g34133 (n_16408, n17982);
  not g34134 (n_16409, n17983);
  and g34135 (n17984, n_16408, n_16409);
  and g34136 (n17985, n_16348, n_16380);
  not g34137 (n_16410, n17985);
  and g34138 (n17986, n17984, n_16410);
  not g34139 (n_16411, n17984);
  and g34140 (n17987, n_16411, n17985);
  not g34141 (n_16412, n17986);
  not g34142 (n_16413, n17987);
  and g34143 (n17988, n_16412, n_16413);
  and g34144 (n17989, \a[46] , \a[63] );
  not g34145 (n_16414, n17891);
  and g34146 (n17990, n_16414, n17989);
  not g34147 (n_16415, n17989);
  and g34148 (n17991, n17891, n_16415);
  not g34149 (n_16416, n17990);
  not g34150 (n_16417, n17991);
  and g34151 (n17992, n_16416, n_16417);
  not g34152 (n_16418, n17992);
  and g34153 (n17993, n17946, n_16418);
  not g34154 (n_16419, n17946);
  and g34155 (n17994, n_16419, n17992);
  not g34156 (n_16420, n17993);
  not g34157 (n_16421, n17994);
  and g34158 (n17995, n_16420, n_16421);
  and g34159 (n17996, n_16324, n_16330);
  not g34160 (n_16422, n17995);
  and g34161 (n17997, n_16422, n17996);
  not g34162 (n_16423, n17996);
  and g34163 (n17998, n17995, n_16423);
  not g34164 (n_16424, n17997);
  not g34165 (n_16425, n17998);
  and g34166 (n17999, n_16424, n_16425);
  and g34167 (n18000, n6325, n9509);
  and g34168 (n18001, n5888, n8905);
  and g34169 (n18002, n6256, n9512);
  not g34170 (n_16426, n18001);
  not g34171 (n_16427, n18002);
  and g34172 (n18003, n_16426, n_16427);
  not g34173 (n_16428, n18000);
  not g34174 (n_16429, n18003);
  and g34175 (n18004, n_16428, n_16429);
  not g34176 (n_16430, n18004);
  and g34177 (n18005, \a[48] , n_16430);
  and g34178 (n18006, \a[61] , n18005);
  and g34179 (n18007, n_16428, n_16430);
  and g34180 (n18008, \a[49] , \a[60] );
  and g34181 (n18009, \a[50] , \a[59] );
  not g34182 (n_16431, n18008);
  not g34183 (n_16432, n18009);
  and g34184 (n18010, n_16431, n_16432);
  not g34185 (n_16433, n18010);
  and g34186 (n18011, n18007, n_16433);
  not g34187 (n_16434, n18006);
  not g34188 (n_16435, n18011);
  and g34189 (n18012, n_16434, n_16435);
  not g34190 (n_16436, n18012);
  and g34191 (n18013, n17927, n_16436);
  not g34192 (n_16437, n17927);
  and g34193 (n18014, n_16437, n18012);
  not g34194 (n_16438, n18013);
  not g34195 (n_16439, n18014);
  and g34196 (n18015, n_16438, n_16439);
  and g34197 (n18016, \a[51] , \a[58] );
  and g34198 (n18017, n7433, n8200);
  and g34199 (n18018, n7232, n7942);
  and g34200 (n18019, n6968, n8436);
  not g34201 (n_16440, n18018);
  not g34202 (n_16441, n18019);
  and g34203 (n18020, n_16440, n_16441);
  not g34204 (n_16442, n18017);
  not g34205 (n_16443, n18020);
  and g34206 (n18021, n_16442, n_16443);
  not g34207 (n_16444, n18021);
  and g34208 (n18022, n18016, n_16444);
  and g34209 (n18023, n_16442, n_16444);
  and g34210 (n18024, \a[52] , \a[57] );
  not g34211 (n_16445, n13288);
  not g34212 (n_16446, n18024);
  and g34213 (n18025, n_16445, n_16446);
  not g34214 (n_16447, n18025);
  and g34215 (n18026, n18023, n_16447);
  not g34216 (n_16448, n18022);
  not g34217 (n_16449, n18026);
  and g34218 (n18027, n_16448, n_16449);
  not g34219 (n_16450, n18015);
  not g34220 (n_16451, n18027);
  and g34221 (n18028, n_16450, n_16451);
  and g34222 (n18029, n18015, n18027);
  not g34223 (n_16452, n18028);
  not g34224 (n_16453, n18029);
  and g34225 (n18030, n_16452, n_16453);
  and g34226 (n18031, n17999, n18030);
  not g34227 (n_16454, n17999);
  not g34228 (n_16455, n18030);
  and g34229 (n18032, n_16454, n_16455);
  not g34230 (n_16456, n18032);
  and g34231 (n18033, n17988, n_16456);
  not g34232 (n_16457, n18031);
  and g34233 (n18034, n_16457, n18033);
  not g34234 (n_16458, n18034);
  and g34235 (n18035, n17988, n_16458);
  and g34236 (n18036, n_16456, n_16458);
  and g34237 (n18037, n_16457, n18036);
  not g34238 (n_16459, n18035);
  not g34239 (n_16460, n18037);
  and g34240 (n18038, n_16459, n_16460);
  and g34241 (n18039, n_16336, n_16381);
  not g34242 (n_16461, n18038);
  not g34243 (n_16462, n18039);
  and g34244 (n18040, n_16461, n_16462);
  and g34245 (n18041, n18038, n18039);
  not g34246 (n_16463, n18040);
  not g34247 (n_16464, n18041);
  and g34248 (n18042, n_16463, n_16464);
  not g34249 (n_16465, n17967);
  not g34250 (n_16466, n18042);
  and g34251 (n18043, n_16465, n_16466);
  and g34252 (n18044, n17967, n18042);
  or g34253 (\asquared[110] , n18043, n18044);
  and g34254 (n18046, n_16465, n_16464);
  not g34255 (n_16467, n18046);
  and g34256 (n18047, n_16463, n_16467);
  and g34257 (n18048, n_16412, n_16458);
  and g34258 (n18049, n18007, n18023);
  not g34259 (n_16468, n18007);
  not g34260 (n_16469, n18023);
  and g34261 (n18050, n_16468, n_16469);
  not g34262 (n_16470, n18049);
  not g34263 (n_16471, n18050);
  and g34264 (n18051, n_16470, n_16471);
  and g34265 (n18052, n6564, n9509);
  and g34266 (n18053, n8905, n9934);
  and g34267 (n18054, n6325, n9512);
  not g34268 (n_16472, n18053);
  not g34269 (n_16473, n18054);
  and g34270 (n18055, n_16472, n_16473);
  not g34271 (n_16474, n18052);
  not g34272 (n_16475, n18055);
  and g34273 (n18056, n_16474, n_16475);
  not g34274 (n_16476, n18056);
  and g34275 (n18057, \a[61] , n_16476);
  and g34276 (n18058, \a[49] , n18057);
  and g34277 (n18059, n_16474, n_16476);
  and g34278 (n18060, \a[50] , \a[60] );
  and g34279 (n18061, \a[51] , \a[59] );
  not g34280 (n_16477, n18060);
  not g34281 (n_16478, n18061);
  and g34282 (n18062, n_16477, n_16478);
  not g34283 (n_16479, n18062);
  and g34284 (n18063, n18059, n_16479);
  not g34285 (n_16480, n18058);
  not g34286 (n_16481, n18063);
  and g34287 (n18064, n_16480, n_16481);
  not g34288 (n_16482, n18064);
  and g34289 (n18065, n18051, n_16482);
  not g34290 (n_16483, n18065);
  and g34291 (n18066, n18051, n_16483);
  and g34292 (n18067, n_16482, n_16483);
  not g34293 (n_16484, n18066);
  not g34294 (n_16485, n18067);
  and g34295 (n18068, n_16484, n_16485);
  and g34296 (n18069, n_16437, n_16436);
  not g34297 (n_16486, n18069);
  and g34298 (n18070, n_16452, n_16486);
  and g34299 (n18071, n18068, n18070);
  not g34300 (n_16487, n18068);
  not g34301 (n_16488, n18070);
  and g34302 (n18072, n_16487, n_16488);
  not g34303 (n_16489, n18071);
  not g34304 (n_16490, n18072);
  and g34305 (n18073, n_16489, n_16490);
  and g34306 (n18074, n_16402, n_16409);
  not g34307 (n_16491, n18073);
  and g34308 (n18075, n_16491, n18074);
  not g34309 (n_16492, n18074);
  and g34310 (n18076, n18073, n_16492);
  not g34311 (n_16493, n18075);
  not g34312 (n_16494, n18076);
  and g34313 (n18077, n_16493, n_16494);
  and g34314 (n18078, n7699, n8200);
  and g34315 (n18079, n7433, n8436);
  and g34316 (n18080, \a[54] , \a[58] );
  and g34317 (n18081, n17892, n18080);
  not g34318 (n_16495, n18079);
  not g34319 (n_16496, n18081);
  and g34320 (n18082, n_16495, n_16496);
  not g34321 (n_16497, n18078);
  not g34322 (n_16498, n18082);
  and g34323 (n18083, n_16497, n_16498);
  not g34324 (n_16499, n18083);
  and g34325 (n18084, \a[58] , n_16499);
  and g34326 (n18085, \a[52] , n18084);
  and g34327 (n18086, n_16497, n_16499);
  and g34328 (n18087, \a[53] , \a[57] );
  not g34329 (n_16500, n7421);
  not g34330 (n_16501, n18087);
  and g34331 (n18088, n_16500, n_16501);
  not g34332 (n_16502, n18088);
  and g34333 (n18089, n18086, n_16502);
  not g34334 (n_16503, n18085);
  not g34335 (n_16504, n18089);
  and g34336 (n18090, n_16503, n_16504);
  and g34337 (n18091, n6252, n9792);
  and g34338 (n18092, \a[47] , \a[63] );
  not g34339 (n_16505, n16400);
  not g34340 (n_16506, n18092);
  and g34341 (n18093, n_16505, n_16506);
  not g34342 (n_16507, n18091);
  not g34343 (n_16508, n18093);
  and g34344 (n18094, n_16507, n_16508);
  not g34345 (n_16509, n17972);
  and g34346 (n18095, n_16509, n18094);
  not g34347 (n_16510, n18094);
  and g34348 (n18096, n17972, n_16510);
  not g34349 (n_16511, n18095);
  not g34350 (n_16512, n18096);
  and g34351 (n18097, n_16511, n_16512);
  not g34352 (n_16513, n18090);
  and g34353 (n18098, n_16513, n18097);
  not g34354 (n_16514, n18098);
  and g34355 (n18099, n18097, n_16514);
  and g34356 (n18100, n_16513, n_16514);
  not g34357 (n_16515, n18099);
  not g34358 (n_16516, n18100);
  and g34359 (n18101, n_16515, n_16516);
  and g34360 (n18102, n_16416, n_16421);
  and g34361 (n18103, n18101, n18102);
  not g34362 (n_16517, n18101);
  not g34363 (n_16518, n18102);
  and g34364 (n18104, n_16517, n_16518);
  not g34365 (n_16519, n18103);
  not g34366 (n_16520, n18104);
  and g34367 (n18105, n_16519, n_16520);
  and g34368 (n18106, n_16425, n_16457);
  not g34369 (n_16521, n18106);
  and g34370 (n18107, n18105, n_16521);
  not g34371 (n_16522, n18107);
  and g34372 (n18108, n18105, n_16522);
  and g34373 (n18109, n_16521, n_16522);
  not g34374 (n_16523, n18108);
  not g34375 (n_16524, n18109);
  and g34376 (n18110, n_16523, n_16524);
  not g34377 (n_16525, n18110);
  and g34378 (n18111, n18077, n_16525);
  not g34379 (n_16526, n18077);
  and g34380 (n18112, n_16526, n_16524);
  and g34381 (n18113, n_16523, n18112);
  not g34382 (n_16527, n18111);
  not g34383 (n_16528, n18113);
  and g34384 (n18114, n_16527, n_16528);
  not g34385 (n_16529, n18114);
  and g34386 (n18115, n18048, n_16529);
  not g34387 (n_16530, n18048);
  and g34388 (n18116, n_16530, n18114);
  not g34389 (n_16531, n18115);
  not g34390 (n_16532, n18116);
  and g34391 (n18117, n_16531, n_16532);
  not g34392 (n_16533, n18117);
  and g34393 (n18118, n18047, n_16533);
  not g34394 (n_16534, n18047);
  and g34395 (n18119, n_16534, n_16531);
  and g34396 (n18120, n_16532, n18119);
  not g34397 (n_16535, n18118);
  not g34398 (n_16536, n18120);
  and g34399 (\asquared[111] , n_16535, n_16536);
  not g34400 (n_16537, n18119);
  and g34401 (n18122, n_16532, n_16537);
  and g34402 (n18123, n_16522, n_16527);
  and g34403 (n18124, n18059, n18086);
  not g34404 (n_16538, n18059);
  not g34405 (n_16539, n18086);
  and g34406 (n18125, n_16538, n_16539);
  not g34407 (n_16540, n18124);
  not g34408 (n_16541, n18125);
  and g34409 (n18126, n_16540, n_16541);
  and g34410 (n18127, n_16507, n_16511);
  not g34411 (n_16542, n18126);
  and g34412 (n18128, n_16542, n18127);
  not g34413 (n_16543, n18127);
  and g34414 (n18129, n18126, n_16543);
  not g34415 (n_16544, n18128);
  not g34416 (n_16545, n18129);
  and g34417 (n18130, n_16544, n_16545);
  and g34418 (n18131, n_16471, n_16483);
  not g34419 (n_16546, n18130);
  and g34420 (n18132, n_16546, n18131);
  not g34421 (n_16547, n18131);
  and g34422 (n18133, n18130, n_16547);
  not g34423 (n_16548, n18132);
  not g34424 (n_16549, n18133);
  and g34425 (n18134, n_16548, n_16549);
  and g34426 (n18135, n_16514, n_16520);
  not g34427 (n_16550, n18134);
  and g34428 (n18136, n_16550, n18135);
  not g34429 (n_16551, n18135);
  and g34430 (n18137, n18134, n_16551);
  not g34431 (n_16552, n18136);
  not g34432 (n_16553, n18137);
  and g34433 (n18138, n_16552, n_16553);
  and g34434 (n18139, n6564, n9512);
  and g34435 (n18140, n11634, n17009);
  and g34436 (n18141, n5888, n9909);
  not g34437 (n_16554, n18140);
  not g34438 (n_16555, n18141);
  and g34439 (n18142, n_16554, n_16555);
  not g34440 (n_16556, n18139);
  not g34441 (n_16557, n18142);
  and g34442 (n18143, n_16556, n_16557);
  not g34443 (n_16558, n18143);
  and g34444 (n18144, n_16556, n_16558);
  and g34445 (n18145, \a[50] , \a[61] );
  and g34446 (n18146, \a[51] , \a[60] );
  not g34447 (n_16559, n18145);
  not g34448 (n_16560, n18146);
  and g34449 (n18147, n_16559, n_16560);
  not g34450 (n_16561, n18147);
  and g34451 (n18148, n18144, n_16561);
  and g34452 (n18149, \a[63] , n_16558);
  and g34453 (n18150, \a[48] , n18149);
  not g34454 (n_16562, n18148);
  not g34455 (n_16563, n18150);
  and g34456 (n18151, n_16562, n_16563);
  and g34457 (n18152, \a[56] , \a[62] );
  and g34458 (n18153, \a[49] , n18152);
  not g34459 (n_16564, n18153);
  and g34460 (n18154, n9161, n_16564);
  not g34461 (n_16565, n18154);
  and g34462 (n18155, n9161, n_16565);
  and g34463 (n18156, n_16564, n_16565);
  not g34464 (n_16566, \a[56] );
  not g34465 (n_16567, n16677);
  and g34466 (n18157, n_16566, n_16567);
  not g34467 (n_16568, n18157);
  and g34468 (n18158, n18156, n_16568);
  not g34469 (n_16569, n18155);
  not g34470 (n_16570, n18158);
  and g34471 (n18159, n_16569, n_16570);
  not g34472 (n_16571, n18151);
  not g34473 (n_16572, n18159);
  and g34474 (n18160, n_16571, n_16572);
  not g34475 (n_16573, n18160);
  and g34476 (n18161, n_16571, n_16573);
  and g34477 (n18162, n_16572, n_16573);
  not g34478 (n_16574, n18161);
  not g34479 (n_16575, n18162);
  and g34480 (n18163, n_16574, n_16575);
  and g34481 (n18164, n7699, n8436);
  and g34482 (n18165, n8985, n10905);
  and g34483 (n18166, n7433, n8987);
  not g34484 (n_16576, n18165);
  not g34485 (n_16577, n18166);
  and g34486 (n18167, n_16576, n_16577);
  not g34487 (n_16578, n18164);
  not g34488 (n_16579, n18167);
  and g34489 (n18168, n_16578, n_16579);
  not g34490 (n_16580, n18168);
  and g34491 (n18169, \a[59] , n_16580);
  and g34492 (n18170, \a[52] , n18169);
  and g34493 (n18171, \a[53] , \a[58] );
  not g34494 (n_16581, n13730);
  not g34495 (n_16582, n18171);
  and g34496 (n18172, n_16581, n_16582);
  and g34497 (n18173, n_16578, n_16580);
  not g34498 (n_16583, n18172);
  and g34499 (n18174, n_16583, n18173);
  not g34500 (n_16584, n18170);
  not g34501 (n_16585, n18174);
  and g34502 (n18175, n_16584, n_16585);
  not g34503 (n_16586, n18163);
  not g34504 (n_16587, n18175);
  and g34505 (n18176, n_16586, n_16587);
  not g34506 (n_16588, n18176);
  and g34507 (n18177, n_16586, n_16588);
  and g34508 (n18178, n_16587, n_16588);
  not g34509 (n_16589, n18177);
  not g34510 (n_16590, n18178);
  and g34511 (n18179, n_16589, n_16590);
  and g34512 (n18180, n_16490, n_16494);
  and g34513 (n18181, n18179, n18180);
  not g34514 (n_16591, n18179);
  not g34515 (n_16592, n18180);
  and g34516 (n18182, n_16591, n_16592);
  not g34517 (n_16593, n18181);
  not g34518 (n_16594, n18182);
  and g34519 (n18183, n_16593, n_16594);
  and g34520 (n18184, n18138, n18183);
  not g34521 (n_16595, n18138);
  not g34522 (n_16596, n18183);
  and g34523 (n18185, n_16595, n_16596);
  not g34524 (n_16597, n18184);
  not g34525 (n_16598, n18185);
  and g34526 (n18186, n_16597, n_16598);
  not g34527 (n_16599, n18123);
  and g34528 (n18187, n_16599, n18186);
  not g34529 (n_16600, n18186);
  and g34530 (n18188, n18123, n_16600);
  not g34531 (n_16601, n18187);
  not g34532 (n_16602, n18188);
  and g34533 (n18189, n_16601, n_16602);
  not g34534 (n_16603, n18122);
  not g34535 (n_16604, n18189);
  and g34536 (n18190, n_16603, n_16604);
  and g34537 (n18191, n18122, n18189);
  or g34538 (\asquared[112] , n18190, n18191);
  and g34539 (n18193, n_16603, n_16602);
  not g34540 (n_16605, n18193);
  and g34541 (n18194, n_16601, n_16605);
  and g34542 (n18195, n_16594, n_16597);
  and g34543 (n18196, n_16549, n_16553);
  and g34544 (n18197, \a[52] , n11634);
  and g34545 (n18198, \a[51] , n9909);
  not g34546 (n_16606, n18197);
  not g34547 (n_16607, n18198);
  and g34548 (n18199, n_16606, n_16607);
  and g34549 (n18200, n6968, n9512);
  not g34550 (n_16608, n18200);
  and g34551 (n18201, \a[49] , n_16608);
  not g34552 (n_16609, n18199);
  and g34553 (n18202, n_16609, n18201);
  not g34554 (n_16610, n18202);
  and g34555 (n18203, \a[49] , n_16610);
  and g34556 (n18204, \a[63] , n18203);
  and g34557 (n18205, n_16608, n_16610);
  and g34558 (n18206, \a[51] , \a[61] );
  and g34559 (n18207, \a[52] , \a[60] );
  not g34560 (n_16611, n18206);
  not g34561 (n_16612, n18207);
  and g34562 (n18208, n_16611, n_16612);
  not g34563 (n_16613, n18208);
  and g34564 (n18209, n18205, n_16613);
  not g34565 (n_16614, n18204);
  not g34566 (n_16615, n18209);
  and g34567 (n18210, n_16614, n_16615);
  not g34568 (n_16616, n18210);
  and g34569 (n18211, n18144, n_16616);
  not g34570 (n_16617, n18144);
  and g34571 (n18212, n_16617, n18210);
  not g34572 (n_16618, n18211);
  not g34573 (n_16619, n18212);
  and g34574 (n18213, n_16618, n_16619);
  and g34575 (n18214, n7701, n8436);
  and g34576 (n18215, n7699, n8987);
  and g34577 (n18216, \a[55] , \a[59] );
  and g34578 (n18217, n18087, n18216);
  not g34579 (n_16620, n18215);
  not g34580 (n_16621, n18217);
  and g34581 (n18218, n_16620, n_16621);
  not g34582 (n_16622, n18214);
  not g34583 (n_16623, n18218);
  and g34584 (n18219, n_16622, n_16623);
  not g34585 (n_16624, n18219);
  and g34586 (n18220, \a[59] , n_16624);
  and g34587 (n18221, \a[53] , n18220);
  and g34588 (n18222, n_16622, n_16624);
  not g34589 (n_16625, n11718);
  not g34590 (n_16626, n18080);
  and g34591 (n18223, n_16625, n_16626);
  not g34592 (n_16627, n18223);
  and g34593 (n18224, n18222, n_16627);
  not g34594 (n_16628, n18221);
  not g34595 (n_16629, n18224);
  and g34596 (n18225, n_16628, n_16629);
  not g34597 (n_16630, n18213);
  not g34598 (n_16631, n18225);
  and g34599 (n18226, n_16630, n_16631);
  and g34600 (n18227, n18213, n18225);
  not g34601 (n_16632, n18226);
  not g34602 (n_16633, n18227);
  and g34603 (n18228, n_16632, n_16633);
  not g34604 (n_16634, n18228);
  and g34605 (n18229, n18196, n_16634);
  not g34606 (n_16635, n18196);
  and g34607 (n18230, n_16635, n18228);
  not g34608 (n_16636, n18229);
  not g34609 (n_16637, n18230);
  and g34610 (n18231, n_16636, n_16637);
  not g34611 (n_16638, n18156);
  and g34612 (n18232, n16921, n_16638);
  not g34613 (n_16639, n16921);
  and g34614 (n18233, n_16639, n18156);
  not g34615 (n_16640, n18232);
  not g34616 (n_16641, n18233);
  and g34617 (n18234, n_16640, n_16641);
  not g34618 (n_16642, n18234);
  and g34619 (n18235, n18173, n_16642);
  not g34620 (n_16643, n18173);
  and g34621 (n18236, n_16643, n18234);
  not g34622 (n_16644, n18235);
  not g34623 (n_16645, n18236);
  and g34624 (n18237, n_16644, n_16645);
  and g34625 (n18238, n_16541, n_16545);
  and g34626 (n18239, n_16573, n_16588);
  and g34627 (n18240, n18238, n18239);
  not g34628 (n_16646, n18238);
  not g34629 (n_16647, n18239);
  and g34630 (n18241, n_16646, n_16647);
  not g34631 (n_16648, n18240);
  not g34632 (n_16649, n18241);
  and g34633 (n18242, n_16648, n_16649);
  and g34634 (n18243, n18237, n18242);
  not g34635 (n_16650, n18237);
  not g34636 (n_16651, n18242);
  and g34637 (n18244, n_16650, n_16651);
  not g34638 (n_16652, n18243);
  not g34639 (n_16653, n18244);
  and g34640 (n18245, n_16652, n_16653);
  and g34641 (n18246, n18231, n18245);
  not g34642 (n_16654, n18231);
  not g34643 (n_16655, n18245);
  and g34644 (n18247, n_16654, n_16655);
  not g34645 (n_16656, n18246);
  not g34646 (n_16657, n18247);
  and g34647 (n18248, n_16656, n_16657);
  not g34648 (n_16658, n18248);
  and g34649 (n18249, n18195, n_16658);
  not g34650 (n_16659, n18195);
  and g34651 (n18250, n_16659, n18248);
  not g34652 (n_16660, n18249);
  not g34653 (n_16661, n18250);
  and g34654 (n18251, n_16660, n_16661);
  not g34655 (n_16662, n18251);
  and g34656 (n18252, n18194, n_16662);
  not g34657 (n_16663, n18194);
  and g34658 (n18253, n_16663, n_16660);
  and g34659 (n18254, n_16661, n18253);
  not g34660 (n_16664, n18252);
  not g34661 (n_16665, n18254);
  and g34662 (\asquared[113] , n_16664, n_16665);
  not g34663 (n_16666, n18253);
  and g34664 (n18256, n_16661, n_16666);
  and g34665 (n18257, n_16637, n_16656);
  and g34666 (n18258, n7433, n9512);
  not g34667 (n_16667, n18258);
  and g34668 (n18259, \a[60] , n_16667);
  and g34669 (n18260, \a[53] , n18259);
  and g34670 (n18261, \a[52] , n_16667);
  and g34671 (n18262, \a[61] , n18261);
  not g34672 (n_16668, n18260);
  not g34673 (n_16669, n18262);
  and g34674 (n18263, n_16668, n_16669);
  not g34675 (n_16670, n18222);
  not g34676 (n_16671, n18263);
  and g34677 (n18264, n_16670, n_16671);
  not g34678 (n_16672, n18264);
  and g34679 (n18265, n_16670, n_16672);
  and g34680 (n18266, n_16671, n_16672);
  not g34681 (n_16673, n18265);
  not g34682 (n_16674, n18266);
  and g34683 (n18267, n_16673, n_16674);
  and g34684 (n18268, n_16640, n_16645);
  and g34685 (n18269, n18267, n18268);
  not g34686 (n_16675, n18267);
  not g34687 (n_16676, n18268);
  and g34688 (n18270, n_16675, n_16676);
  not g34689 (n_16677, n18269);
  not g34690 (n_16678, n18270);
  and g34691 (n18271, n_16677, n_16678);
  and g34692 (n18272, n_16617, n_16616);
  not g34693 (n_16679, n18272);
  and g34694 (n18273, n_16632, n_16679);
  not g34695 (n_16680, n18271);
  and g34696 (n18274, n_16680, n18273);
  not g34697 (n_16681, n18273);
  and g34698 (n18275, n18271, n_16681);
  not g34699 (n_16682, n18274);
  not g34700 (n_16683, n18275);
  and g34701 (n18276, n_16682, n_16683);
  and g34702 (n18277, n_16649, n_16652);
  and g34703 (n18278, \a[54] , \a[59] );
  not g34704 (n_16684, n16457);
  not g34705 (n_16685, n18278);
  and g34706 (n18279, n_16684, n_16685);
  and g34707 (n18280, n7701, n8987);
  not g34708 (n_16686, n18280);
  not g34711 (n_16687, n18279);
  not g34713 (n_16688, n18283);
  and g34714 (n18284, \a[50] , n_16688);
  and g34715 (n18285, \a[63] , n18284);
  and g34716 (n18286, n_16686, n_16688);
  and g34717 (n18287, n_16687, n18286);
  not g34718 (n_16689, n18285);
  not g34719 (n_16690, n18287);
  and g34720 (n18288, n_16689, n_16690);
  not g34721 (n_16691, n18288);
  and g34722 (n18289, n18205, n_16691);
  not g34723 (n_16692, n18205);
  and g34724 (n18290, n_16692, n18288);
  not g34725 (n_16693, n18289);
  not g34726 (n_16694, n18290);
  and g34727 (n18291, n_16693, n_16694);
  and g34728 (n18292, \a[62] , n14417);
  not g34729 (n_16695, n18292);
  and g34730 (n18293, n8200, n_16695);
  not g34731 (n_16696, n18293);
  and g34732 (n18294, n8200, n_16696);
  and g34733 (n18295, n_16695, n_16696);
  not g34734 (n_16697, \a[57] );
  not g34735 (n_16698, n14081);
  and g34736 (n18296, n_16697, n_16698);
  not g34737 (n_16699, n18296);
  and g34738 (n18297, n18295, n_16699);
  not g34739 (n_16700, n18294);
  not g34740 (n_16701, n18297);
  and g34741 (n18298, n_16700, n_16701);
  not g34742 (n_16702, n18291);
  not g34743 (n_16703, n18298);
  and g34744 (n18299, n_16702, n_16703);
  and g34745 (n18300, n18291, n18298);
  not g34746 (n_16704, n18299);
  not g34747 (n_16705, n18300);
  and g34748 (n18301, n_16704, n_16705);
  not g34749 (n_16706, n18277);
  and g34750 (n18302, n_16706, n18301);
  not g34751 (n_16707, n18301);
  and g34752 (n18303, n18277, n_16707);
  not g34753 (n_16708, n18302);
  not g34754 (n_16709, n18303);
  and g34755 (n18304, n_16708, n_16709);
  not g34756 (n_16710, n18276);
  not g34757 (n_16711, n18304);
  and g34758 (n18305, n_16710, n_16711);
  and g34759 (n18306, n18276, n18304);
  not g34760 (n_16712, n18305);
  not g34761 (n_16713, n18306);
  and g34762 (n18307, n_16712, n_16713);
  not g34763 (n_16714, n18307);
  and g34764 (n18308, n18257, n_16714);
  not g34765 (n_16715, n18257);
  and g34766 (n18309, n_16715, n18307);
  not g34767 (n_16716, n18308);
  not g34768 (n_16717, n18309);
  and g34769 (n18310, n_16716, n_16717);
  not g34770 (n_16718, n18256);
  not g34771 (n_16719, n18310);
  and g34772 (n18311, n_16718, n_16719);
  and g34773 (n18312, n18256, n18310);
  or g34774 (\asquared[114] , n18311, n18312);
  and g34775 (n18314, n_16718, n_16716);
  not g34776 (n_16720, n18314);
  and g34777 (n18315, n_16717, n_16720);
  and g34778 (n18316, n_16708, n_16713);
  and g34779 (n18317, n18286, n18295);
  not g34780 (n_16721, n18286);
  not g34781 (n_16722, n18295);
  and g34782 (n18318, n_16721, n_16722);
  not g34783 (n_16723, n18317);
  not g34784 (n_16724, n18318);
  and g34785 (n18319, n_16723, n_16724);
  and g34786 (n18320, n_16667, n_16672);
  not g34787 (n_16725, n18319);
  and g34788 (n18321, n_16725, n18320);
  not g34789 (n_16726, n18320);
  and g34790 (n18322, n18319, n_16726);
  not g34791 (n_16727, n18321);
  not g34792 (n_16728, n18322);
  and g34793 (n18323, n_16727, n_16728);
  and g34794 (n18324, n_16678, n_16683);
  not g34795 (n_16729, n18323);
  and g34796 (n18325, n_16729, n18324);
  not g34797 (n_16730, n18324);
  and g34798 (n18326, n18323, n_16730);
  not g34799 (n_16731, n18325);
  not g34800 (n_16732, n18326);
  and g34801 (n18327, n_16731, n_16732);
  and g34802 (n18328, \a[52] , \a[62] );
  and g34803 (n18329, \a[53] , \a[61] );
  not g34804 (n_16733, n18328);
  not g34805 (n_16734, n18329);
  and g34806 (n18330, n_16733, n_16734);
  and g34807 (n18331, n7433, n9721);
  and g34808 (n18332, n6968, n9792);
  and g34809 (n18333, n7232, n9909);
  not g34810 (n_16735, n18332);
  not g34811 (n_16736, n18333);
  and g34812 (n18334, n_16735, n_16736);
  not g34813 (n_16737, n18331);
  not g34814 (n_16738, n18334);
  and g34815 (n18335, n_16737, n_16738);
  not g34816 (n_16739, n18335);
  and g34817 (n18336, n_16737, n_16739);
  not g34818 (n_16740, n18330);
  and g34819 (n18337, n_16740, n18336);
  and g34820 (n18338, \a[63] , n_16739);
  and g34821 (n18339, \a[51] , n18338);
  not g34822 (n_16741, n18337);
  not g34823 (n_16742, n18339);
  and g34824 (n18340, n_16741, n_16742);
  and g34825 (n18341, n8987, n9161);
  and g34826 (n18342, n7421, n10089);
  and g34827 (n18343, n7701, n9509);
  not g34828 (n_16743, n18342);
  not g34829 (n_16744, n18343);
  and g34830 (n18344, n_16743, n_16744);
  not g34831 (n_16745, n18341);
  not g34832 (n_16746, n18344);
  and g34833 (n18345, n_16745, n_16746);
  not g34834 (n_16747, n18345);
  and g34835 (n18346, \a[60] , n_16747);
  and g34836 (n18347, \a[54] , n18346);
  and g34837 (n18348, n_16745, n_16747);
  not g34838 (n_16748, n7942);
  not g34839 (n_16749, n18216);
  and g34840 (n18349, n_16748, n_16749);
  not g34841 (n_16750, n18349);
  and g34842 (n18350, n18348, n_16750);
  not g34843 (n_16751, n18347);
  not g34844 (n_16752, n18350);
  and g34845 (n18351, n_16751, n_16752);
  not g34846 (n_16753, n18340);
  not g34847 (n_16754, n18351);
  and g34848 (n18352, n_16753, n_16754);
  not g34849 (n_16755, n18352);
  and g34850 (n18353, n_16753, n_16755);
  and g34851 (n18354, n_16754, n_16755);
  not g34852 (n_16756, n18353);
  not g34853 (n_16757, n18354);
  and g34854 (n18355, n_16756, n_16757);
  and g34855 (n18356, n_16692, n_16691);
  not g34856 (n_16758, n18356);
  and g34857 (n18357, n_16704, n_16758);
  and g34858 (n18358, n18355, n18357);
  not g34859 (n_16759, n18355);
  not g34860 (n_16760, n18357);
  and g34861 (n18359, n_16759, n_16760);
  not g34862 (n_16761, n18358);
  not g34863 (n_16762, n18359);
  and g34864 (n18360, n_16761, n_16762);
  and g34865 (n18361, n18327, n18360);
  not g34866 (n_16763, n18327);
  not g34867 (n_16764, n18360);
  and g34868 (n18362, n_16763, n_16764);
  not g34869 (n_16765, n18361);
  not g34870 (n_16766, n18362);
  and g34871 (n18363, n_16765, n_16766);
  not g34872 (n_16767, n18363);
  and g34873 (n18364, n18316, n_16767);
  not g34874 (n_16768, n18316);
  and g34875 (n18365, n_16768, n18363);
  not g34876 (n_16769, n18364);
  not g34877 (n_16770, n18365);
  and g34878 (n18366, n_16769, n_16770);
  not g34879 (n_16771, n18366);
  and g34880 (n18367, n18315, n_16771);
  not g34881 (n_16772, n18315);
  and g34882 (n18368, n_16772, n_16769);
  and g34883 (n18369, n_16770, n18368);
  not g34884 (n_16773, n18367);
  not g34885 (n_16774, n18369);
  and g34886 (\asquared[115] , n_16773, n_16774);
  not g34887 (n_16775, n18368);
  and g34888 (n18371, n_16770, n_16775);
  and g34889 (n18372, n_16732, n_16765);
  and g34890 (n18373, \a[53] , \a[62] );
  and g34891 (n18374, \a[58] , n18373);
  not g34892 (n_16776, n18374);
  and g34893 (n18375, n8436, n_16776);
  not g34894 (n_16777, n18375);
  and g34895 (n18376, n_16776, n_16777);
  not g34896 (n_16778, \a[58] );
  not g34897 (n_16779, n18373);
  and g34898 (n18377, n_16778, n_16779);
  not g34899 (n_16780, n18377);
  and g34900 (n18378, n18376, n_16780);
  and g34901 (n18379, n8436, n_16777);
  not g34902 (n_16781, n18378);
  not g34903 (n_16782, n18379);
  and g34904 (n18380, n_16781, n_16782);
  and g34905 (n18381, n9161, n9509);
  and g34906 (n18382, n7421, n8905);
  and g34907 (n18383, n7701, n9512);
  not g34908 (n_16783, n18382);
  not g34909 (n_16784, n18383);
  and g34910 (n18384, n_16783, n_16784);
  not g34911 (n_16785, n18381);
  not g34912 (n_16786, n18384);
  and g34913 (n18385, n_16785, n_16786);
  not g34914 (n_16787, n18385);
  and g34915 (n18386, \a[61] , n_16787);
  and g34916 (n18387, \a[54] , n18386);
  and g34917 (n18388, n_16785, n_16787);
  and g34918 (n18389, \a[55] , \a[60] );
  not g34919 (n_16788, n13870);
  not g34920 (n_16789, n18389);
  and g34921 (n18390, n_16788, n_16789);
  not g34922 (n_16790, n18390);
  and g34923 (n18391, n18388, n_16790);
  not g34924 (n_16791, n18387);
  not g34925 (n_16792, n18391);
  and g34926 (n18392, n_16791, n_16792);
  not g34927 (n_16793, n18380);
  not g34928 (n_16794, n18392);
  and g34929 (n18393, n_16793, n_16794);
  not g34930 (n_16795, n18393);
  and g34931 (n18394, n_16793, n_16795);
  and g34932 (n18395, n_16794, n_16795);
  not g34933 (n_16796, n18394);
  not g34934 (n_16797, n18395);
  and g34935 (n18396, n_16796, n_16797);
  and g34936 (n18397, n_16724, n_16728);
  and g34937 (n18398, n18396, n18397);
  not g34938 (n_16798, n18396);
  not g34939 (n_16799, n18397);
  and g34940 (n18399, n_16798, n_16799);
  not g34941 (n_16800, n18398);
  not g34942 (n_16801, n18399);
  and g34943 (n18400, n_16800, n_16801);
  and g34944 (n18401, \a[52] , \a[63] );
  not g34945 (n_16802, n18348);
  and g34946 (n18402, n_16802, n18401);
  not g34947 (n_16803, n18401);
  and g34948 (n18403, n18348, n_16803);
  not g34949 (n_16804, n18402);
  not g34950 (n_16805, n18403);
  and g34951 (n18404, n_16804, n_16805);
  not g34952 (n_16806, n18404);
  and g34953 (n18405, n18336, n_16806);
  not g34954 (n_16807, n18336);
  and g34955 (n18406, n_16807, n18404);
  not g34956 (n_16808, n18405);
  not g34957 (n_16809, n18406);
  and g34958 (n18407, n_16808, n_16809);
  and g34959 (n18408, n_16755, n_16762);
  not g34960 (n_16810, n18407);
  and g34961 (n18409, n_16810, n18408);
  not g34962 (n_16811, n18408);
  and g34963 (n18410, n18407, n_16811);
  not g34964 (n_16812, n18409);
  not g34965 (n_16813, n18410);
  and g34966 (n18411, n_16812, n_16813);
  and g34967 (n18412, n18400, n18411);
  not g34968 (n_16814, n18400);
  not g34969 (n_16815, n18411);
  and g34970 (n18413, n_16814, n_16815);
  not g34971 (n_16816, n18412);
  not g34972 (n_16817, n18413);
  and g34973 (n18414, n_16816, n_16817);
  not g34974 (n_16818, n18372);
  and g34975 (n18415, n_16818, n18414);
  not g34976 (n_16819, n18414);
  and g34977 (n18416, n18372, n_16819);
  not g34978 (n_16820, n18415);
  not g34979 (n_16821, n18416);
  and g34980 (n18417, n_16820, n_16821);
  not g34981 (n_16822, n18371);
  not g34982 (n_16823, n18417);
  and g34983 (n18418, n_16822, n_16823);
  and g34984 (n18419, n18371, n18417);
  or g34985 (\asquared[116] , n18418, n18419);
  and g34986 (n18421, n_16822, n_16821);
  not g34987 (n_16824, n18421);
  and g34988 (n18422, n_16820, n_16824);
  and g34989 (n18423, n_16795, n_16801);
  and g34990 (n18424, n_16804, n_16809);
  and g34991 (n18425, n18423, n18424);
  not g34992 (n_16825, n18423);
  not g34993 (n_16826, n18424);
  and g34994 (n18426, n_16825, n_16826);
  not g34995 (n_16827, n18425);
  not g34996 (n_16828, n18426);
  and g34997 (n18427, n_16827, n_16828);
  and g34998 (n18428, n7699, n9792);
  not g34999 (n_16829, n18428);
  and g35000 (n18429, \a[62] , n_16829);
  and g35001 (n18430, \a[54] , n18429);
  and g35002 (n18431, \a[53] , n_16829);
  and g35003 (n18432, \a[63] , n18431);
  not g35004 (n_16830, n18430);
  not g35005 (n_16831, n18432);
  and g35006 (n18433, n_16830, n_16831);
  not g35007 (n_16832, n18376);
  not g35008 (n_16833, n18433);
  and g35009 (n18434, n_16832, n_16833);
  not g35010 (n_16834, n18434);
  and g35011 (n18435, n_16832, n_16834);
  and g35012 (n18436, n_16833, n_16834);
  not g35013 (n_16835, n18435);
  not g35014 (n_16836, n18436);
  and g35015 (n18437, n_16835, n_16836);
  and g35016 (n18438, n8200, n9509);
  and g35017 (n18439, n8905, n11718);
  and g35018 (n18440, n9161, n9512);
  not g35019 (n_16837, n18439);
  not g35020 (n_16838, n18440);
  and g35021 (n18441, n_16837, n_16838);
  not g35022 (n_16839, n18438);
  not g35023 (n_16840, n18441);
  and g35024 (n18442, n_16839, n_16840);
  not g35025 (n_16841, n18442);
  and g35026 (n18443, \a[55] , n_16841);
  and g35027 (n18444, \a[61] , n18443);
  and g35028 (n18445, n_16839, n_16841);
  and g35029 (n18446, \a[56] , \a[60] );
  not g35030 (n_16842, n8985);
  not g35031 (n_16843, n18446);
  and g35032 (n18447, n_16842, n_16843);
  not g35033 (n_16844, n18447);
  and g35034 (n18448, n18445, n_16844);
  not g35035 (n_16845, n18444);
  not g35036 (n_16846, n18448);
  and g35037 (n18449, n_16845, n_16846);
  not g35038 (n_16847, n18388);
  not g35039 (n_16848, n18449);
  and g35040 (n18450, n_16847, n_16848);
  not g35041 (n_16849, n18450);
  and g35042 (n18451, n_16847, n_16849);
  and g35043 (n18452, n_16848, n_16849);
  not g35044 (n_16850, n18451);
  not g35045 (n_16851, n18452);
  and g35046 (n18453, n_16850, n_16851);
  not g35047 (n_16852, n18437);
  not g35048 (n_16853, n18453);
  and g35049 (n18454, n_16852, n_16853);
  and g35050 (n18455, n18437, n_16851);
  and g35051 (n18456, n_16850, n18455);
  not g35052 (n_16854, n18454);
  not g35053 (n_16855, n18456);
  and g35054 (n18457, n_16854, n_16855);
  and g35055 (n18458, n18427, n18457);
  not g35056 (n_16856, n18427);
  not g35057 (n_16857, n18457);
  and g35058 (n18459, n_16856, n_16857);
  not g35059 (n_16858, n18458);
  not g35060 (n_16859, n18459);
  and g35061 (n18460, n_16858, n_16859);
  and g35062 (n18461, n_16813, n_16816);
  not g35063 (n_16860, n18460);
  and g35064 (n18462, n_16860, n18461);
  not g35065 (n_16861, n18461);
  and g35066 (n18463, n18460, n_16861);
  not g35067 (n_16862, n18462);
  not g35068 (n_16863, n18463);
  and g35069 (n18464, n_16862, n_16863);
  not g35070 (n_16864, n18464);
  and g35071 (n18465, n18422, n_16864);
  not g35072 (n_16865, n18422);
  and g35073 (n18466, n_16865, n_16862);
  and g35074 (n18467, n_16863, n18466);
  not g35075 (n_16866, n18465);
  not g35076 (n_16867, n18467);
  and g35077 (\asquared[117] , n_16866, n_16867);
  not g35078 (n_16868, n18466);
  and g35079 (n18469, n_16863, n_16868);
  and g35080 (n18470, n_16828, n_16858);
  and g35081 (n18471, n_16829, n_16834);
  and g35082 (n18472, n18445, n18471);
  not g35083 (n_16869, n18445);
  not g35084 (n_16870, n18471);
  and g35085 (n18473, n_16869, n_16870);
  not g35086 (n_16871, n18472);
  not g35087 (n_16872, n18473);
  and g35088 (n18474, n_16871, n_16872);
  and g35089 (n18475, n8200, n9512);
  and g35090 (n18476, n11634, n13730);
  and g35091 (n18477, n7421, n9909);
  not g35092 (n_16873, n18476);
  not g35093 (n_16874, n18477);
  and g35094 (n18478, n_16873, n_16874);
  not g35095 (n_16875, n18475);
  not g35096 (n_16876, n18478);
  and g35097 (n18479, n_16875, n_16876);
  not g35098 (n_16877, n18479);
  and g35099 (n18480, \a[63] , n_16877);
  and g35100 (n18481, \a[54] , n18480);
  and g35101 (n18482, \a[56] , \a[61] );
  not g35102 (n_16878, n13212);
  not g35103 (n_16879, n18482);
  and g35104 (n18483, n_16878, n_16879);
  and g35105 (n18484, n_16875, n_16877);
  not g35106 (n_16880, n18483);
  and g35107 (n18485, n_16880, n18484);
  not g35108 (n_16881, n18481);
  not g35109 (n_16882, n18485);
  and g35110 (n18486, n_16881, n_16882);
  not g35111 (n_16883, n18486);
  and g35112 (n18487, n18474, n_16883);
  not g35113 (n_16884, n18487);
  and g35114 (n18488, n18474, n_16884);
  and g35115 (n18489, n_16883, n_16884);
  not g35116 (n_16885, n18488);
  not g35117 (n_16886, n18489);
  and g35118 (n18490, n_16885, n_16886);
  and g35119 (n18491, n_16849, n_16854);
  and g35120 (n18492, \a[55] , n16295);
  not g35121 (n_16887, n18492);
  and g35122 (n18493, n8987, n_16887);
  not g35123 (n_16888, n18493);
  and g35124 (n18494, n8987, n_16888);
  and g35125 (n18495, n_16887, n_16888);
  and g35126 (n18496, \a[55] , \a[62] );
  not g35127 (n_16889, \a[59] );
  not g35128 (n_16890, n18496);
  and g35129 (n18497, n_16889, n_16890);
  not g35130 (n_16891, n18497);
  and g35131 (n18498, n18495, n_16891);
  not g35132 (n_16892, n18494);
  not g35133 (n_16893, n18498);
  and g35134 (n18499, n_16892, n_16893);
  not g35135 (n_16894, n18491);
  not g35136 (n_16895, n18499);
  and g35137 (n18500, n_16894, n_16895);
  not g35138 (n_16896, n18500);
  and g35139 (n18501, n_16894, n_16896);
  and g35140 (n18502, n_16895, n_16896);
  not g35141 (n_16897, n18501);
  not g35142 (n_16898, n18502);
  and g35143 (n18503, n_16897, n_16898);
  not g35144 (n_16899, n18490);
  and g35145 (n18504, n_16899, n18503);
  not g35146 (n_16900, n18503);
  and g35147 (n18505, n18490, n_16900);
  not g35148 (n_16901, n18504);
  not g35149 (n_16902, n18505);
  and g35150 (n18506, n_16901, n_16902);
  not g35151 (n_16903, n18470);
  not g35152 (n_16904, n18506);
  and g35153 (n18507, n_16903, n_16904);
  and g35154 (n18508, n18470, n18506);
  not g35155 (n_16905, n18507);
  not g35156 (n_16906, n18508);
  and g35157 (n18509, n_16905, n_16906);
  not g35158 (n_16907, n18469);
  not g35159 (n_16908, n18509);
  and g35160 (n18510, n_16907, n_16908);
  and g35161 (n18511, n18469, n18509);
  or g35162 (\asquared[118] , n18510, n18511);
  and g35163 (n18513, \a[55] , \a[63] );
  not g35164 (n_16909, n18495);
  and g35165 (n18514, n_16909, n18513);
  not g35166 (n_16910, n18513);
  and g35167 (n18515, n18495, n_16910);
  not g35168 (n_16911, n18514);
  not g35169 (n_16912, n18515);
  and g35170 (n18516, n_16911, n_16912);
  not g35171 (n_16913, n18516);
  and g35172 (n18517, n18484, n_16913);
  not g35173 (n_16914, n18484);
  and g35174 (n18518, n_16914, n18516);
  not g35175 (n_16915, n18517);
  not g35176 (n_16916, n18518);
  and g35177 (n18519, n_16915, n_16916);
  and g35178 (n18520, n_16872, n_16884);
  and g35179 (n18521, n8436, n9512);
  and g35180 (n18522, n10089, n18152);
  and g35181 (n18523, n8200, n9721);
  not g35182 (n_16917, n18522);
  not g35183 (n_16918, n18523);
  and g35184 (n18524, n_16917, n_16918);
  not g35185 (n_16919, n18521);
  not g35186 (n_16920, n18524);
  and g35187 (n18525, n_16919, n_16920);
  not g35188 (n_16921, n18525);
  and g35189 (n18526, n18152, n_16921);
  and g35190 (n18527, n_16919, n_16921);
  and g35191 (n18528, \a[57] , \a[61] );
  not g35192 (n_16922, n10089);
  not g35193 (n_16923, n18528);
  and g35194 (n18529, n_16922, n_16923);
  not g35195 (n_16924, n18529);
  and g35196 (n18530, n18527, n_16924);
  not g35197 (n_16925, n18526);
  not g35198 (n_16926, n18530);
  and g35199 (n18531, n_16925, n_16926);
  not g35200 (n_16927, n18520);
  not g35201 (n_16928, n18531);
  and g35202 (n18532, n_16927, n_16928);
  not g35203 (n_16929, n18532);
  and g35204 (n18533, n_16927, n_16929);
  and g35205 (n18534, n_16928, n_16929);
  not g35206 (n_16930, n18533);
  not g35207 (n_16931, n18534);
  and g35208 (n18535, n_16930, n_16931);
  not g35209 (n_16932, n18519);
  and g35210 (n18536, n_16932, n18535);
  not g35211 (n_16933, n18535);
  and g35212 (n18537, n18519, n_16933);
  not g35213 (n_16934, n18536);
  not g35214 (n_16935, n18537);
  and g35215 (n18538, n_16934, n_16935);
  and g35216 (n18539, n_16899, n_16900);
  not g35217 (n_16936, n18539);
  and g35218 (n18540, n_16896, n_16936);
  not g35219 (n_16937, n18538);
  and g35220 (n18541, n_16937, n18540);
  not g35221 (n_16938, n18540);
  and g35222 (n18542, n18538, n_16938);
  not g35223 (n_16939, n18541);
  not g35224 (n_16940, n18542);
  and g35225 (n18543, n_16939, n_16940);
  and g35226 (n18544, n_16907, n_16906);
  not g35227 (n_16941, n18544);
  and g35228 (n18545, n_16905, n_16941);
  not g35229 (n_16942, n18543);
  and g35230 (n18546, n_16942, n18545);
  not g35231 (n_16943, n18545);
  and g35232 (n18547, n18543, n_16943);
  not g35233 (n_16944, n18546);
  not g35234 (n_16945, n18547);
  and g35235 (\asquared[119] , n_16944, n_16945);
  and g35236 (n18549, n7942, n9909);
  not g35237 (n_16946, n18549);
  and g35238 (n18550, \a[61] , n_16946);
  and g35239 (n18551, \a[58] , n18550);
  and g35240 (n18552, \a[56] , n_16946);
  and g35241 (n18553, \a[63] , n18552);
  not g35242 (n_16947, n18551);
  not g35243 (n_16948, n18553);
  and g35244 (n18554, n_16947, n_16948);
  not g35245 (n_16949, n18527);
  not g35246 (n_16950, n18554);
  and g35247 (n18555, n_16949, n_16950);
  not g35248 (n_16951, n18555);
  and g35249 (n18556, n_16949, n_16951);
  and g35250 (n18557, n_16950, n_16951);
  not g35251 (n_16952, n18556);
  not g35252 (n_16953, n18557);
  and g35253 (n18558, n_16952, n_16953);
  and g35254 (n18559, \a[57] , n9085);
  not g35255 (n_16954, n18559);
  and g35256 (n18560, n9509, n_16954);
  not g35257 (n_16955, n18560);
  and g35258 (n18561, n9509, n_16955);
  and g35259 (n18562, n_16954, n_16955);
  and g35260 (n18563, \a[57] , \a[62] );
  not g35261 (n_16956, \a[60] );
  not g35262 (n_16957, n18563);
  and g35263 (n18564, n_16956, n_16957);
  not g35264 (n_16958, n18564);
  and g35265 (n18565, n18562, n_16958);
  not g35266 (n_16959, n18561);
  not g35267 (n_16960, n18565);
  and g35268 (n18566, n_16959, n_16960);
  not g35269 (n_16961, n18558);
  not g35270 (n_16962, n18566);
  and g35271 (n18567, n_16961, n_16962);
  not g35272 (n_16963, n18567);
  and g35273 (n18568, n_16961, n_16963);
  and g35274 (n18569, n_16962, n_16963);
  not g35275 (n_16964, n18568);
  not g35276 (n_16965, n18569);
  and g35277 (n18570, n_16964, n_16965);
  and g35278 (n18571, n_16911, n_16916);
  and g35279 (n18572, n18570, n18571);
  not g35280 (n_16966, n18570);
  not g35281 (n_16967, n18571);
  and g35282 (n18573, n_16966, n_16967);
  not g35283 (n_16968, n18572);
  not g35284 (n_16969, n18573);
  and g35285 (n18574, n_16968, n_16969);
  and g35286 (n18575, n_16929, n_16935);
  not g35287 (n_16970, n18575);
  and g35288 (n18576, n18574, n_16970);
  not g35289 (n_16971, n18574);
  and g35290 (n18577, n_16971, n18575);
  not g35291 (n_16972, n18576);
  not g35292 (n_16973, n18577);
  and g35293 (n18578, n_16972, n_16973);
  and g35294 (n18579, n_16939, n_16943);
  not g35295 (n_16974, n18579);
  and g35296 (n18580, n_16940, n_16974);
  not g35297 (n_16975, n18578);
  and g35298 (n18581, n_16975, n18580);
  not g35299 (n_16976, n18580);
  and g35300 (n18582, n18578, n_16976);
  not g35301 (n_16977, n18581);
  not g35302 (n_16978, n18582);
  and g35303 (\asquared[120] , n_16977, n_16978);
  and g35304 (n18584, n_16973, n_16976);
  not g35305 (n_16979, n18584);
  and g35306 (n18585, n_16972, n_16979);
  and g35307 (n18586, n_16963, n_16969);
  and g35308 (n18587, n_16946, n_16951);
  and g35309 (n18588, n18562, n18587);
  not g35310 (n_16980, n18562);
  not g35311 (n_16981, n18587);
  and g35312 (n18589, n_16980, n_16981);
  not g35313 (n_16982, n18588);
  not g35314 (n_16983, n18589);
  and g35315 (n18590, n_16982, n_16983);
  and g35316 (n18591, n8987, n9721);
  and g35317 (n18592, n8985, n9909);
  and g35318 (n18593, n8436, n9792);
  not g35319 (n_16984, n18592);
  not g35320 (n_16985, n18593);
  and g35321 (n18594, n_16984, n_16985);
  not g35322 (n_16986, n18591);
  not g35323 (n_16987, n18594);
  and g35324 (n18595, n_16986, n_16987);
  not g35325 (n_16988, n18595);
  and g35326 (n18596, \a[63] , n_16988);
  and g35327 (n18597, \a[57] , n18596);
  and g35328 (n18598, n_16986, n_16988);
  and g35329 (n18599, \a[58] , \a[62] );
  not g35330 (n_16989, n8905);
  not g35331 (n_16990, n18599);
  and g35332 (n18600, n_16989, n_16990);
  not g35333 (n_16991, n18600);
  and g35334 (n18601, n18598, n_16991);
  not g35335 (n_16992, n18597);
  not g35336 (n_16993, n18601);
  and g35337 (n18602, n_16992, n_16993);
  not g35338 (n_16994, n18602);
  and g35339 (n18603, n18590, n_16994);
  not g35340 (n_16995, n18590);
  and g35341 (n18604, n_16995, n18602);
  not g35342 (n_16996, n18603);
  not g35343 (n_16997, n18604);
  and g35344 (n18605, n_16996, n_16997);
  not g35345 (n_16998, n18605);
  and g35346 (n18606, n18586, n_16998);
  not g35347 (n_16999, n18586);
  and g35348 (n18607, n_16999, n18605);
  not g35349 (n_17000, n18606);
  not g35350 (n_17001, n18607);
  and g35351 (n18608, n_17000, n_17001);
  not g35352 (n_17002, n18608);
  and g35353 (n18609, n18585, n_17002);
  not g35354 (n_17003, n18585);
  and g35355 (n18610, n_17003, n_17000);
  and g35356 (n18611, n_17001, n18610);
  not g35357 (n_17004, n18609);
  not g35358 (n_17005, n18611);
  and g35359 (\asquared[121] , n_17004, n_17005);
  and g35360 (n18613, n_16956, \a[61] );
  not g35361 (n_17006, n16295);
  not g35362 (n_17007, n18613);
  and g35363 (n18614, n_17006, n_17007);
  and g35364 (n18615, n16295, n18613);
  not g35365 (n_17008, n18614);
  not g35366 (n_17009, n18615);
  and g35367 (n18616, n_17008, n_17009);
  not g35368 (n_17010, n18598);
  and g35369 (n18617, n17799, n_17010);
  not g35370 (n_17011, n17799);
  and g35371 (n18618, n_17011, n18598);
  not g35372 (n_17012, n18617);
  not g35373 (n_17013, n18618);
  and g35374 (n18619, n_17012, n_17013);
  not g35375 (n_17014, n18616);
  not g35376 (n_17015, n18619);
  and g35377 (n18620, n_17014, n_17015);
  and g35378 (n18621, n18616, n18619);
  not g35379 (n_17016, n18620);
  not g35380 (n_17017, n18621);
  and g35381 (n18622, n_17016, n_17017);
  and g35382 (n18623, n_16983, n_16996);
  not g35383 (n_17018, n18622);
  and g35384 (n18624, n_17018, n18623);
  not g35385 (n_17019, n18623);
  and g35386 (n18625, n18622, n_17019);
  not g35387 (n_17020, n18624);
  not g35388 (n_17021, n18625);
  and g35389 (n18626, n_17020, n_17021);
  not g35390 (n_17022, n18610);
  and g35391 (n18627, n_17001, n_17022);
  not g35392 (n_17023, n18626);
  and g35393 (n18628, n_17023, n18627);
  not g35394 (n_17024, n18627);
  and g35395 (n18629, n18626, n_17024);
  not g35396 (n_17025, n18628);
  not g35397 (n_17026, n18629);
  and g35398 (\asquared[122] , n_17025, n_17026);
  and g35399 (n18631, n_17020, n_17024);
  not g35400 (n_17027, n18631);
  and g35401 (n18632, n_17021, n_17027);
  not g35402 (n_17028, n9085);
  not g35403 (n_17029, n17802);
  and g35404 (n18633, n_17028, n_17029);
  and g35405 (n18634, n9509, n9792);
  not g35406 (n_17030, n9512);
  and g35407 (n18635, n_17030, n_17009);
  not g35408 (n_17031, n18634);
  not g35409 (n_17032, n18635);
  and g35410 (n18636, n_17031, n_17032);
  not g35411 (n_17033, n18633);
  and g35412 (n18637, n_17033, n18636);
  not g35413 (n_17034, n18637);
  and g35414 (n18638, n_17031, n_17034);
  and g35415 (n18639, n_17033, n18638);
  and g35416 (n18640, n_17032, n_17034);
  not g35417 (n_17035, n18639);
  not g35418 (n_17036, n18640);
  and g35419 (n18641, n_17035, n_17036);
  and g35420 (n18642, n_17012, n_17017);
  and g35421 (n18643, n18641, n18642);
  not g35422 (n_17037, n18641);
  not g35423 (n_17038, n18642);
  and g35424 (n18644, n_17037, n_17038);
  not g35425 (n_17039, n18643);
  not g35426 (n_17040, n18644);
  and g35427 (n18645, n_17039, n_17040);
  not g35428 (n_17041, n18645);
  and g35429 (n18646, n18632, n_17041);
  not g35430 (n_17042, n18632);
  and g35431 (n18647, n_17042, n_17039);
  and g35432 (n18648, n_17040, n18647);
  not g35433 (n_17043, n18646);
  not g35434 (n_17044, n18648);
  and g35435 (\asquared[123] , n_17043, n_17044);
  not g35436 (n_17045, \a[61] );
  and g35437 (n18650, n_17045, \a[62] );
  not g35438 (n_17046, n11634);
  not g35439 (n_17047, n18650);
  and g35440 (n18651, n_17046, n_17047);
  and g35441 (n18652, n11634, n18650);
  not g35442 (n_17048, n18651);
  not g35443 (n_17049, n18652);
  and g35444 (n18653, n_17048, n_17049);
  not g35445 (n_17050, n18653);
  and g35446 (n18654, n18638, n_17050);
  not g35447 (n_17051, n18638);
  and g35448 (n18655, n_17051, n18653);
  not g35449 (n_17052, n18654);
  not g35450 (n_17053, n18655);
  and g35451 (n18656, n_17052, n_17053);
  not g35452 (n_17054, n18647);
  and g35453 (n18657, n_17040, n_17054);
  not g35454 (n_17055, n18656);
  and g35455 (n18658, n_17055, n18657);
  not g35456 (n_17056, n18657);
  and g35457 (n18659, n18656, n_17056);
  not g35458 (n_17057, n18658);
  not g35459 (n_17058, n18659);
  and g35460 (\asquared[124] , n_17057, n_17058);
  and g35461 (n18661, n_17052, n_17056);
  not g35462 (n_17059, n18661);
  and g35463 (n18662, n_17053, n_17059);
  and g35464 (n18663, \a[62] , n9909);
  not g35465 (n_17060, n9721);
  not g35466 (n_17061, n9909);
  and g35467 (n18664, n_17060, n_17061);
  and g35468 (n18665, n_17049, n18664);
  not g35469 (n_17062, n18663);
  not g35470 (n_17063, n18665);
  and g35471 (n18666, n_17062, n_17063);
  not g35472 (n_17064, n18662);
  and g35473 (n18667, n_17064, n18666);
  not g35474 (n_17065, n18666);
  and g35475 (n18668, n18662, n_17065);
  not g35476 (n_17066, n18667);
  not g35477 (n_17067, n18668);
  and g35478 (\asquared[125] , n_17066, n_17067);
  not g35479 (n_17068, \a[62] );
  and g35480 (n18670, n_17068, \a[63] );
  and g35481 (n18671, n_17064, n_17063);
  not g35482 (n_17069, n18671);
  and g35483 (n18672, n_17062, n_17069);
  not g35484 (n_17070, n18670);
  and g35485 (n18673, n_17070, n18672);
  not g35486 (n_17071, n18672);
  and g35487 (n18674, n18670, n_17071);
  not g35488 (n_17072, n18673);
  not g35489 (n_17073, n18674);
  and g35490 (\asquared[126] , n_17072, n_17073);
  and g35491 (n18676, \a[63] , n_17071);
  or g35492 (\asquared[127] , n9792, n18676);
  and g35493 (n667, n_428, \a[13] , \a[2] , n_427);
  and g35494 (n1254, n_963, \a[22] , \a[0] , n_961);
  and g35495 (n1610, n_1287, \a[20] , \a[5] , n_1286);
  and g35496 (n1802, n_1461, \a[22] , \a[5] , n_1460);
  and g35497 (n1908, n_1563, \a[20] , \a[8] , n_1562);
  and g35498 (n2091, n_1725, \a[12] , \a[17] , n_1724);
  and g35499 (n2200, n_1827, \a[13] , \a[17] , n_1826);
  and g35500 (n2321, n_1933, \a[25] , \a[6] , n_1932);
  and g35501 (n2519, n_2108, \a[14] , \a[18] , n_2107);
  and g35502 (n2457, n_2059, \a[9] , \a[23] , n_2058);
  and g35503 (n2655, n_2244, \a[26] , \a[7] , n_2243);
  and g35504 (n2754, n_2336, \a[32] , \a[2] , n_2335);
  and g35505 (n2955, n_2518, \a[31] , \a[4] , n_2517);
  and g35506 (n2939, n_2506, \a[28] , \a[7] , n_2505);
  and g35507 (n3085, n_2638, \a[34] , \a[2] , n_2637);
  and g35508 (n3323, n_2851, \a[16] , \a[21] , n_2850);
  and g35509 (n3283, n_2820, \a[29] , \a[8] , n_2819);
  and g35510 (n3547, n_3055, \a[35] , \a[3] , n_3054);
  and g35511 (n3642, n_3152, \a[17] , \a[22] , n_3151);
  and g35512 (n3653, n_3159, \a[31] , \a[8] , n_3158);
  and g35513 (n3860, n_3347, \a[37] , \a[3] , n_3346);
  and g35514 (n4002, n_3487, \a[38] , \a[3] , n_3486);
  and g35515 (n4041, n_3517, \a[33] , \a[8] , n_3516);
  and g35516 (n4444, n_3878, \a[41] , \a[2] , n_3877);
  and g35517 (n4428, n_3866, \a[9] , \a[34] , n_3865);
  and g35518 (n4617, n_4032, \a[39] , \a[5] , n_4031);
  and g35519 (n4537, n_3970, \a[41] , \a[3] , n_3969);
  and g35520 (n4844, n_4247, \a[10] , \a[35] , n_4246);
  and g35521 (n4963, n_4356, \a[44] , \a[2] , n_4355);
  and g35522 (n5332, n_4693, \a[10] , \a[37] , n_4692);
  and g35523 (n5625, n_4961, \a[13] , \a[36] , n_4960);
  and g35524 (n5635, n_4968, \a[11] , \a[38] , n_4967);
  and g35525 (n5670, n_4995, \a[22] , \a[27] , n_4994);
  and g35526 (n6102, \a[17] , n_5398, \a[34] , n_5401);
  and g35527 (n6201, n_5482, \a[11] , \a[40] , n_5481);
  and g35528 (n6329, n_5608, \a[19] , \a[33] , n_5607);
  and g35529 (n6474, n_5744, \a[15] , \a[37] , n_5743);
  and g35530 (n6646, n_5893, \a[53] , \a[0] , n_5891);
  and g35531 (n6693, n_5934, \a[11] , \a[42] , n_5933);
  and g35532 (n6578, n_5836, \a[49] , \a[4] , n_5835);
  and g35533 (n7218, n_6426, \a[16] , \a[39] , n_6425);
  and g35534 (n7151, n_6367, \a[50] , \a[5] , n_6366);
  and g35535 (n7202, n_6414, \a[12] , \a[43] , n_6413);
  and g35536 (n7067, n_6290, \a[52] , \a[3] , n_6289);
  and g35537 (n7540, n_6718, \a[21] , \a[35] , n_6717);
  and g35538 (n7735, n_6894, \a[15] , \a[42] , n_6893);
  and g35539 (n7719, n_6882, \a[52] , \a[5] , n_6881);
  and g35540 (n7762, n_6916, \a[12] , \a[45] , n_6915);
  and g35541 (n8087, n_7217, \a[55] , \a[3] , n_7216);
  and g35542 (n7996, n_7135, \a[18] , \a[40] , n_7134);
  and g35543 (n7962, n_7108, \a[53] , \a[5] , n_7107);
  and g35544 (n8187, n_7307, \a[51] , \a[8] , n_7306);
  and g35545 (n8889, n_7952, \a[13] , \a[48] , n_7951);
  and g35546 (n8925, n_7979, \a[55] , \a[6] , n_7978);
  and g35547 (n8752, n_7818, \a[23] , \a[38] , n_7817);
  and g35548 (n8694, n_7771, \a[19] , \a[42] , n_7770);
  and g35549 (n9165, n_8182, \a[20] , \a[42] , n_8181);
  and g35550 (n9533, n_8525, \a[58] , \a[5] , n_8524);
  and g35551 (n9469, n_8477, \a[23] , \a[40] , n_8476);
  and g35552 (n9480, n_8484, \a[14] , \a[49] , n_8483);
  and g35553 (n9670, n_8656, \a[26] , \a[38] , n_8655);
  and g35554 (n10078, n_9034, \a[57] , \a[8] , n_9033);
  and g35555 (n10039, n_9000, \a[36] , \a[29] , n_8999);
  and g35556 (n10340, n_9278, \a[10] , \a[56] , n_9277);
  and g35557 (n10356, n_9290, \a[18] , \a[48] , n_9289);
  and g35558 (n10367, n_9297, \a[14] , \a[52] , n_9296);
  and g35559 (n10477, n_9398, \a[63] , \a[4] , n_9397);
  and g35560 (n10848, n_9755, \a[21] , \a[47] , n_9754);
  and g35561 (n10921, \a[48] , n_9811, \a[20] , n_9814);
  and g35562 (n11144, n_10016, \a[14] , \a[55] , n_10015);
  and g35563 (n11107, n_9986, \a[63] , \a[6] , n_9985);
  and g35564 (n11303, n_10175, \a[28] , \a[42] , n_10174);
  and g35565 (n11336, n_10201, \a[22] , \a[48] , n_10200);
  and g35566 (n11697, n_10540, \a[23] , \a[48] , n_10539);
  and g35567 (n11592, n_10448, \a[22] , \a[49] , n_10447);
  and g35568 (n11917, n_10744, \a[12] , \a[60] , n_10743);
  and g35569 (n11861, n_10700, \a[40] , \a[32] , n_10699);
  and g35570 (n12166, n_10976, \a[17] , \a[56] , n_10975);
  and g35571 (n12107, n_10929, \a[23] , \a[50] , n_10928);
  and g35572 (n12204, n_11012, \a[25] , \a[48] , n_11011);
  and g35573 (n12347, \a[11] , n_11141, \a[63] , n_11140);
  and g35574 (n12551, n_11339, \a[30] , \a[45] , n_11338);
  and g35575 (n12673, n_11445, \a[41] , \a[34] , n_11444);
  and g35576 (n12883, n_11640, \a[18] , \a[58] , n_11639);
  and g35577 (n12912, \a[13] , n_11660, \a[63] , n_11659);
  and g35578 (n13163, n_11892, \a[16] , \a[61] , n_11891);
  and g35579 (n13135, n_11870, \a[34] , \a[43] , n_11869);
  and g35580 (n13371, n_12087, \a[23] , \a[55] , n_12086);
  and g35581 (n13265, n_11980, \a[20] , \a[58] , n_11979);
  and g35582 (n13548, n_12253, \a[28] , \a[51] , n_12252);
  and g35583 (n13448, n_12161, \a[16] , \a[63] , n_12160);
  and g35584 (n13660, n_12352, \a[47] , \a[33] , n_12351);
  and g35585 (n14138, n_12792, \a[26] , \a[56] , n_12791);
  and g35586 (n14383, n_13034, \a[29] , \a[54] , n_13033);
  and g35587 (n14538, n_13170, \a[51] , \a[33] , n_13169);
  and g35588 (n14692, n_13312, \a[35] , \a[50] , n_13311);
  and g35589 (n14989, n_13589, \a[30] , \a[56] , n_13588);
  and g35590 (n14921, \a[23] , n_13530, \a[63] , n_13529);
  and g35591 (n15172, n_13761, \a[32] , \a[55] , n_13760);
  and g35592 (n15122, n_13720, \a[40] , \a[47] , n_13719);
  and g35593 (n15261, n_13838, \a[57] , \a[31] , n_13837);
  and g35594 (n15294, n_13865, \a[59] , \a[29] , n_13864);
  and g35595 (n15551, \a[26] , n_14105, \a[63] , n_14104);
  and g35596 (n15419, n_13986, \a[41] , \a[48] , n_13985);
  and g35597 (n15834, n_14374, \a[28] , \a[63] , n_14373);
  and g35598 (n15846, n_14381, \a[35] , \a[56] , n_14380);
  and g35599 (n16040, \a[32] , \a[60] , n_14558, n_14559);
  and g35600 (n16254, n_14768, \a[58] , \a[36] , n_14767);
  and g35601 (n16450, n_14951, \a[41] , \a[54] , n_14950);
  and g35602 (n16414, \a[39] , \a[56] , n_14919, n_14920);
  and g35603 (n16691, n_15179, \a[40] , \a[57] , n_15178);
  and g35604 (n16820, n_15303, \a[53] , \a[45] , n_15302);
  and g35605 (n17169, n_15634, \a[63] , \a[38] , n_15633);
  and g35606 (n17404, n_15850, \a[60] , \a[43] , n_15849);
  and g35607 (n18283, n_16687, \a[63] , \a[50] , n_16686);
endmodule

