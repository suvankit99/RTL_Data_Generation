
module Priority(\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] ,
     \A[7] , \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14]
     , \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] ,
     \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] ,
     \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] ,
     \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] ,
     \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] ,
     \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
     \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
     \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] ,
     \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] ,
     \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] ,
     \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] ,
     \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] ,
     \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] , \A[105]
     , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] , \A[111] ,
     \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
     \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
     \A[124] , \A[125] , \A[126] , \A[127] , \P[0] , \P[1] , \P[2] ,
     \P[3] , \P[4] , \P[5] , \P[6] , F);
  input \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
       \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] ,
       \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] ,
       \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] ,
       \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] ,
       \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] ,
       \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] ,
       \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
       \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
       \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] ,
       \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] ,
       \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] ,
       \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] ,
       \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] ,
       \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] ,
       \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
       \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
       \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] ,
       \A[123] , \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
       \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] ,
       \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] ,
       \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] ,
       \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] ,
       \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] ,
       \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] ,
       \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
       \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
       \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] ,
       \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] ,
       \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] ,
       \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] ,
       \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] ,
       \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] ,
       \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
       \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
       \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] ,
       \A[123] , \A[124] , \A[125] , \A[126] , \A[127] ;
  wire \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire n137, n138, n139, n140, n141, n142, n143, n144;
  wire n145, n146, n147, n148, n149, n150, n151, n152;
  wire n153, n154, n155, n156, n157, n158, n159, n160;
  wire n161, n162, n163, n164, n165, n166, n167, n168;
  wire n169, n170, n171, n172, n173, n174, n175, n176;
  wire n177, n178, n179, n180, n181, n182, n183, n184;
  wire n185, n186, n187, n188, n189, n190, n191, n192;
  wire n193, n194, n195, n196, n197, n198, n199, n200;
  wire n201, n202, n203, n204, n205, n206, n207, n208;
  wire n209, n210, n211, n212, n213, n214, n215, n216;
  wire n217, n218, n219, n220, n221, n222, n223, n224;
  wire n225, n226, n227, n228, n229, n230, n231, n232;
  wire n233, n234, n235, n236, n237, n238, n239, n240;
  wire n241, n242, n243, n244, n245, n246, n247, n248;
  wire n249, n250, n251, n252, n253, n254, n255, n256;
  wire n257, n258, n259, n260, n261, n262, n263, n264;
  wire n265, n266, n267, n268, n269, n270, n271, n272;
  wire n273, n274, n275, n276, n277, n278, n279, n280;
  wire n281, n282, n283, n284, n285, n286, n287, n288;
  wire n289, n290, n291, n292, n293, n294, n295, n296;
  wire n297, n298, n299, n300, n301, n302, n303, n304;
  wire n305, n306, n307, n308, n309, n310, n311, n312;
  wire n313, n314, n315, n316, n317, n318, n319, n320;
  wire n321, n322, n323, n324, n325, n326, n327, n328;
  wire n329, n330, n331, n332, n333, n334, n335, n336;
  wire n337, n338, n339, n340, n341, n342, n343, n344;
  wire n345, n346, n347, n348, n349, n350, n351, n352;
  wire n353, n354, n355, n356, n357, n358, n359, n360;
  wire n361, n362, n363, n364, n365, n366, n367, n368;
  wire n369, n370, n371, n372, n373, n374, n375, n376;
  wire n377, n378, n379, n380, n381, n382, n383, n384;
  wire n385, n386, n387, n388, n389, n390, n391, n392;
  wire n393, n394, n395, n396, n397, n398, n399, n400;
  wire n401, n402, n403, n404, n405, n406, n407, n408;
  wire n409, n410, n411, n412, n413, n414, n415, n416;
  wire n417, n418, n419, n420, n421, n422, n423, n424;
  wire n425, n426, n427, n428, n429, n430, n431, n432;
  wire n433, n434, n435, n436, n437, n438, n439, n440;
  wire n441, n442, n443, n444, n445, n446, n447, n448;
  wire n449, n450, n451, n452, n453, n454, n455, n456;
  wire n457, n458, n459, n460, n461, n462, n463, n464;
  wire n465, n466, n467, n468, n469, n470, n471, n472;
  wire n473, n474, n475, n476, n477, n478, n479, n480;
  wire n481, n482, n483, n484, n485, n486, n487, n488;
  wire n489, n490, n491, n492, n493, n494, n495, n496;
  wire n497, n498, n499, n500, n501, n502, n503, n504;
  wire n505, n506, n507, n508, n509, n510, n512, n513;
  wire n514, n515, n516, n517, n518, n519, n520, n521;
  wire n522, n523, n524, n525, n526, n527, n528, n529;
  wire n530, n531, n532, n533, n534, n535, n536, n537;
  wire n538, n539, n540, n541, n542, n543, n544, n545;
  wire n546, n547, n548, n549, n550, n551, n552, n553;
  wire n554, n555, n556, n557, n558, n559, n560, n561;
  wire n562, n563, n564, n565, n566, n567, n568, n569;
  wire n570, n571, n572, n573, n574, n575, n576, n577;
  wire n578, n579, n580, n581, n582, n583, n584, n585;
  wire n586, n587, n588, n589, n590, n591, n592, n593;
  wire n594, n595, n596, n597, n598, n599, n600, n601;
  wire n602, n603, n604, n605, n606, n607, n608, n609;
  wire n610, n611, n612, n613, n614, n615, n616, n617;
  wire n618, n619, n620, n621, n622, n623, n624, n625;
  wire n626, n627, n628, n629, n630, n631, n632, n633;
  wire n634, n635, n636, n637, n638, n639, n640, n641;
  wire n642, n643, n644, n645, n646, n647, n648, n649;
  wire n650, n651, n652, n653, n654, n655, n656, n657;
  wire n658, n659, n660, n661, n662, n663, n664, n665;
  wire n666, n667, n668, n669, n670, n671, n672, n673;
  wire n674, n675, n676, n677, n678, n679, n680, n681;
  wire n682, n683, n684, n685, n686, n687, n688, n689;
  wire n690, n691, n692, n693, n694, n695, n696, n697;
  wire n698, n699, n700, n701, n702, n703, n704, n705;
  wire n706, n707, n708, n709, n710, n711, n712, n713;
  wire n714, n715, n716, n717, n718, n719, n720, n721;
  wire n722, n723, n724, n725, n726, n727, n728, n729;
  wire n730, n731, n732, n733, n734, n735, n736, n737;
  wire n738, n739, n740, n741, n742, n743, n744, n745;
  wire n746, n747, n748, n749, n750, n751, n752, n753;
  wire n754, n755, n756, n757, n758, n760, n761, n762;
  wire n763, n764, n765, n766, n767, n768, n769, n770;
  wire n771, n772, n773, n774, n775, n776, n777, n778;
  wire n779, n780, n781, n782, n783, n784, n785, n786;
  wire n787, n788, n789, n790, n791, n792, n793, n794;
  wire n795, n796, n797, n798, n799, n800, n801, n802;
  wire n803, n804, n805, n806, n807, n808, n809, n810;
  wire n811, n812, n813, n814, n815, n816, n817, n818;
  wire n819, n820, n821, n822, n823, n824, n825, n826;
  wire n827, n828, n829, n830, n831, n832, n833, n834;
  wire n835, n836, n837, n838, n839, n840, n841, n842;
  wire n843, n844, n845, n846, n847, n848, n849, n850;
  wire n851, n852, n853, n854, n855, n856, n857, n858;
  wire n859, n860, n861, n862, n863, n864, n865, n866;
  wire n867, n868, n869, n870, n871, n872, n873, n874;
  wire n875, n876, n877, n878, n879, n880, n881, n882;
  wire n883, n884, n885, n886, n887, n888, n889, n890;
  wire n891, n892, n893, n894, n895, n896, n897, n898;
  wire n899, n900, n901, n902, n903, n904, n905, n906;
  wire n907, n908, n910, n913, n917, n918, n919, n925;
  wire n926, n927, n928, n929, n930, n931, n935, n936;
  wire n937, n938, n942, n943, n944, n945, n949, n950;
  wire n951, n952, n956, n957, n958, n959, n963, n964;
  wire n965, n966, n970, n971, n972, n973, n977, n978;
  wire n979, n980, n984, n985, n986, n987, n991, n992;
  wire n993, n994, n998, n999, n1000, n1001, n1005, n1006;
  wire n1007, n1009, n1014, n1022, n1023, n1024, n1038, n1039;
  wire n1040, n1041, n1042, n1043, n1044, n1052, n1053, n1054;
  wire n1055, n1063, n1064, n1065, n1066, n1074, n1075, n1076;
  wire n1078, n1087, n1103, n1104, n_2, n_5, n_6, n_7;
  wire n_8, n_10, n_11, n_13, n_14, n_15, n_16, n_17;
  wire n_18, n_20, n_21, n_23, n_24, n_25, n_26, n_27;
  wire n_28, n_30, n_31, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_40, n_41, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_50, n_51, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_60, n_61, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_70, n_71, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_80, n_81, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_90, n_91, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_100, n_101, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_110, n_111, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_120, n_121, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_130, n_131, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_140, n_141, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_150, n_151, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_160, n_161, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_170, n_171, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_180, n_181, n_183, n_184, n_185, n_186, n_187;
  wire n_188, n_190, n_191, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_200, n_201, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_210, n_211, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_220, n_221, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_230, n_231, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_240, n_241, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_250, n_251, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_260, n_261, n_263, n_264, n_265, n_266, n_267;
  wire n_268, n_270, n_271, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_280, n_281, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_290, n_291, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_300, n_301, n_303, n_304, n_305, n_306, n_307;
  wire n_308, n_310, n_311, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_320, n_321, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_330, n_331, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_340, n_341, n_343, n_344, n_345, n_346, n_347;
  wire n_348, n_350, n_351, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_360, n_361, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_370, n_371, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_380, n_381, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_390, n_391, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_400, n_401, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_410, n_411, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_420, n_421, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_430, n_431, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_440, n_441, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_450, n_451, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_460, n_461, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_470, n_471, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_480, n_481, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_490, n_491, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_500, n_501, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  wire n_518, n_520, n_521, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_530, n_531, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_540, n_541, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_550, n_551, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_560, n_561, n_563, n_564, n_565, n_566, n_567;
  wire n_568, n_570, n_571, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_580, n_581, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_590, n_591, n_593, n_594, n_595, n_596, n_597;
  wire n_598, n_600, n_601, n_603, n_604, n_605, n_606, n_607;
  wire n_608, n_610, n_611, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_621, n_622, n_623, n_624, n_625, n_626, n_627;
  wire n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659;
  wire n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  wire n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787;
  wire n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811;
  wire n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819;
  wire n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835;
  wire n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843;
  wire n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867;
  wire n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875;
  wire n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883;
  wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
  wire n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899;
  wire n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907;
  wire n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915;
  wire n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923;
  wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931;
  wire n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939;
  wire n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947;
  wire n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955;
  wire n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963;
  wire n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971;
  wire n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979;
  wire n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003;
  wire n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011;
  wire n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019;
  wire n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043;
  wire n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088;
  wire n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096;
  wire n_1097, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1106;
  wire n_1108, n_1109, n_1110, n_1111, n_1113, n_1114, n_1115, n_1116;
  not g1 (n_2, \A[125] );
  and g2 (n137, n_2, \A[127] );
  and g3 (n138, \A[126] , \A[127] );
  not g4 (n_5, n138);
  and g5 (n139, \A[126] , n_5);
  not g6 (n_6, n139);
  and g7 (n140, \A[125] , n_6);
  not g8 (n_7, n137);
  not g9 (n_8, n140);
  and g10 (n141, n_7, n_8);
  not g11 (n_10, \A[123] );
  not g12 (n_11, n141);
  and g13 (n142, n_10, n_11);
  not g14 (n_13, \A[124] );
  and g15 (n143, n_13, n_6);
  and g16 (n144, \A[124] , n_11);
  not g17 (n_14, n143);
  not g18 (n_15, n144);
  and g19 (n145, n_14, n_15);
  not g20 (n_16, n145);
  and g21 (n146, \A[123] , n_16);
  not g22 (n_17, n142);
  not g23 (n_18, n146);
  and g24 (n147, n_17, n_18);
  not g25 (n_20, \A[121] );
  not g26 (n_21, n147);
  and g27 (n148, n_20, n_21);
  not g28 (n_23, \A[122] );
  and g29 (n149, n_23, n_16);
  and g30 (n150, \A[122] , n_21);
  not g31 (n_24, n149);
  not g32 (n_25, n150);
  and g33 (n151, n_24, n_25);
  not g34 (n_26, n151);
  and g35 (n152, \A[121] , n_26);
  not g36 (n_27, n148);
  not g37 (n_28, n152);
  and g38 (n153, n_27, n_28);
  not g39 (n_30, \A[119] );
  not g40 (n_31, n153);
  and g41 (n154, n_30, n_31);
  not g42 (n_33, \A[120] );
  and g43 (n155, n_33, n_26);
  and g44 (n156, \A[120] , n_31);
  not g45 (n_34, n155);
  not g46 (n_35, n156);
  and g47 (n157, n_34, n_35);
  not g48 (n_36, n157);
  and g49 (n158, \A[119] , n_36);
  not g50 (n_37, n154);
  not g51 (n_38, n158);
  and g52 (n159, n_37, n_38);
  not g53 (n_40, \A[117] );
  not g54 (n_41, n159);
  and g55 (n160, n_40, n_41);
  not g56 (n_43, \A[118] );
  and g57 (n161, n_43, n_36);
  and g58 (n162, \A[118] , n_41);
  not g59 (n_44, n161);
  not g60 (n_45, n162);
  and g61 (n163, n_44, n_45);
  not g62 (n_46, n163);
  and g63 (n164, \A[117] , n_46);
  not g64 (n_47, n160);
  not g65 (n_48, n164);
  and g66 (n165, n_47, n_48);
  not g67 (n_50, \A[115] );
  not g68 (n_51, n165);
  and g69 (n166, n_50, n_51);
  not g70 (n_53, \A[116] );
  and g71 (n167, n_53, n_46);
  and g72 (n168, \A[116] , n_51);
  not g73 (n_54, n167);
  not g74 (n_55, n168);
  and g75 (n169, n_54, n_55);
  not g76 (n_56, n169);
  and g77 (n170, \A[115] , n_56);
  not g78 (n_57, n166);
  not g79 (n_58, n170);
  and g80 (n171, n_57, n_58);
  not g81 (n_60, \A[113] );
  not g82 (n_61, n171);
  and g83 (n172, n_60, n_61);
  not g84 (n_63, \A[114] );
  and g85 (n173, n_63, n_56);
  and g86 (n174, \A[114] , n_61);
  not g87 (n_64, n173);
  not g88 (n_65, n174);
  and g89 (n175, n_64, n_65);
  not g90 (n_66, n175);
  and g91 (n176, \A[113] , n_66);
  not g92 (n_67, n172);
  not g93 (n_68, n176);
  and g94 (n177, n_67, n_68);
  not g95 (n_70, \A[111] );
  not g96 (n_71, n177);
  and g97 (n178, n_70, n_71);
  not g98 (n_73, \A[112] );
  and g99 (n179, n_73, n_66);
  and g100 (n180, \A[112] , n_71);
  not g101 (n_74, n179);
  not g102 (n_75, n180);
  and g103 (n181, n_74, n_75);
  not g104 (n_76, n181);
  and g105 (n182, \A[111] , n_76);
  not g106 (n_77, n178);
  not g107 (n_78, n182);
  and g108 (n183, n_77, n_78);
  not g109 (n_80, \A[109] );
  not g110 (n_81, n183);
  and g111 (n184, n_80, n_81);
  not g112 (n_83, \A[110] );
  and g113 (n185, n_83, n_76);
  and g114 (n186, \A[110] , n_81);
  not g115 (n_84, n185);
  not g116 (n_85, n186);
  and g117 (n187, n_84, n_85);
  not g118 (n_86, n187);
  and g119 (n188, \A[109] , n_86);
  not g120 (n_87, n184);
  not g121 (n_88, n188);
  and g122 (n189, n_87, n_88);
  not g123 (n_90, \A[107] );
  not g124 (n_91, n189);
  and g125 (n190, n_90, n_91);
  not g126 (n_93, \A[108] );
  and g127 (n191, n_93, n_86);
  and g128 (n192, \A[108] , n_91);
  not g129 (n_94, n191);
  not g130 (n_95, n192);
  and g131 (n193, n_94, n_95);
  not g132 (n_96, n193);
  and g133 (n194, \A[107] , n_96);
  not g134 (n_97, n190);
  not g135 (n_98, n194);
  and g136 (n195, n_97, n_98);
  not g137 (n_100, \A[105] );
  not g138 (n_101, n195);
  and g139 (n196, n_100, n_101);
  not g140 (n_103, \A[106] );
  and g141 (n197, n_103, n_96);
  and g142 (n198, \A[106] , n_101);
  not g143 (n_104, n197);
  not g144 (n_105, n198);
  and g145 (n199, n_104, n_105);
  not g146 (n_106, n199);
  and g147 (n200, \A[105] , n_106);
  not g148 (n_107, n196);
  not g149 (n_108, n200);
  and g150 (n201, n_107, n_108);
  not g151 (n_110, \A[103] );
  not g152 (n_111, n201);
  and g153 (n202, n_110, n_111);
  not g154 (n_113, \A[104] );
  and g155 (n203, n_113, n_106);
  and g156 (n204, \A[104] , n_111);
  not g157 (n_114, n203);
  not g158 (n_115, n204);
  and g159 (n205, n_114, n_115);
  not g160 (n_116, n205);
  and g161 (n206, \A[103] , n_116);
  not g162 (n_117, n202);
  not g163 (n_118, n206);
  and g164 (n207, n_117, n_118);
  not g165 (n_120, \A[101] );
  not g166 (n_121, n207);
  and g167 (n208, n_120, n_121);
  not g168 (n_123, \A[102] );
  and g169 (n209, n_123, n_116);
  and g170 (n210, \A[102] , n_121);
  not g171 (n_124, n209);
  not g172 (n_125, n210);
  and g173 (n211, n_124, n_125);
  not g174 (n_126, n211);
  and g175 (n212, \A[101] , n_126);
  not g176 (n_127, n208);
  not g177 (n_128, n212);
  and g178 (n213, n_127, n_128);
  not g179 (n_130, \A[99] );
  not g180 (n_131, n213);
  and g181 (n214, n_130, n_131);
  not g182 (n_133, \A[100] );
  and g183 (n215, n_133, n_126);
  and g184 (n216, \A[100] , n_131);
  not g185 (n_134, n215);
  not g186 (n_135, n216);
  and g187 (n217, n_134, n_135);
  not g188 (n_136, n217);
  and g189 (n218, \A[99] , n_136);
  not g190 (n_137, n214);
  not g191 (n_138, n218);
  and g192 (n219, n_137, n_138);
  not g193 (n_140, \A[97] );
  not g194 (n_141, n219);
  and g195 (n220, n_140, n_141);
  not g196 (n_143, \A[98] );
  and g197 (n221, n_143, n_136);
  and g198 (n222, \A[98] , n_141);
  not g199 (n_144, n221);
  not g200 (n_145, n222);
  and g201 (n223, n_144, n_145);
  not g202 (n_146, n223);
  and g203 (n224, \A[97] , n_146);
  not g204 (n_147, n220);
  not g205 (n_148, n224);
  and g206 (n225, n_147, n_148);
  not g207 (n_150, \A[95] );
  not g208 (n_151, n225);
  and g209 (n226, n_150, n_151);
  not g210 (n_153, \A[96] );
  and g211 (n227, n_153, n_146);
  and g212 (n228, \A[96] , n_151);
  not g213 (n_154, n227);
  not g214 (n_155, n228);
  and g215 (n229, n_154, n_155);
  not g216 (n_156, n229);
  and g217 (n230, \A[95] , n_156);
  not g218 (n_157, n226);
  not g219 (n_158, n230);
  and g220 (n231, n_157, n_158);
  not g221 (n_160, \A[93] );
  not g222 (n_161, n231);
  and g223 (n232, n_160, n_161);
  not g224 (n_163, \A[94] );
  and g225 (n233, n_163, n_156);
  and g226 (n234, \A[94] , n_161);
  not g227 (n_164, n233);
  not g228 (n_165, n234);
  and g229 (n235, n_164, n_165);
  not g230 (n_166, n235);
  and g231 (n236, \A[93] , n_166);
  not g232 (n_167, n232);
  not g233 (n_168, n236);
  and g234 (n237, n_167, n_168);
  not g235 (n_170, \A[91] );
  not g236 (n_171, n237);
  and g237 (n238, n_170, n_171);
  not g238 (n_173, \A[92] );
  and g239 (n239, n_173, n_166);
  and g240 (n240, \A[92] , n_171);
  not g241 (n_174, n239);
  not g242 (n_175, n240);
  and g243 (n241, n_174, n_175);
  not g244 (n_176, n241);
  and g245 (n242, \A[91] , n_176);
  not g246 (n_177, n238);
  not g247 (n_178, n242);
  and g248 (n243, n_177, n_178);
  not g249 (n_180, \A[89] );
  not g250 (n_181, n243);
  and g251 (n244, n_180, n_181);
  not g252 (n_183, \A[90] );
  and g253 (n245, n_183, n_176);
  and g254 (n246, \A[90] , n_181);
  not g255 (n_184, n245);
  not g256 (n_185, n246);
  and g257 (n247, n_184, n_185);
  not g258 (n_186, n247);
  and g259 (n248, \A[89] , n_186);
  not g260 (n_187, n244);
  not g261 (n_188, n248);
  and g262 (n249, n_187, n_188);
  not g263 (n_190, \A[87] );
  not g264 (n_191, n249);
  and g265 (n250, n_190, n_191);
  not g266 (n_193, \A[88] );
  and g267 (n251, n_193, n_186);
  and g268 (n252, \A[88] , n_191);
  not g269 (n_194, n251);
  not g270 (n_195, n252);
  and g271 (n253, n_194, n_195);
  not g272 (n_196, n253);
  and g273 (n254, \A[87] , n_196);
  not g274 (n_197, n250);
  not g275 (n_198, n254);
  and g276 (n255, n_197, n_198);
  not g277 (n_200, \A[85] );
  not g278 (n_201, n255);
  and g279 (n256, n_200, n_201);
  not g280 (n_203, \A[86] );
  and g281 (n257, n_203, n_196);
  and g282 (n258, \A[86] , n_201);
  not g283 (n_204, n257);
  not g284 (n_205, n258);
  and g285 (n259, n_204, n_205);
  not g286 (n_206, n259);
  and g287 (n260, \A[85] , n_206);
  not g288 (n_207, n256);
  not g289 (n_208, n260);
  and g290 (n261, n_207, n_208);
  not g291 (n_210, \A[83] );
  not g292 (n_211, n261);
  and g293 (n262, n_210, n_211);
  not g294 (n_213, \A[84] );
  and g295 (n263, n_213, n_206);
  and g296 (n264, \A[84] , n_211);
  not g297 (n_214, n263);
  not g298 (n_215, n264);
  and g299 (n265, n_214, n_215);
  not g300 (n_216, n265);
  and g301 (n266, \A[83] , n_216);
  not g302 (n_217, n262);
  not g303 (n_218, n266);
  and g304 (n267, n_217, n_218);
  not g305 (n_220, \A[81] );
  not g306 (n_221, n267);
  and g307 (n268, n_220, n_221);
  not g308 (n_223, \A[82] );
  and g309 (n269, n_223, n_216);
  and g310 (n270, \A[82] , n_221);
  not g311 (n_224, n269);
  not g312 (n_225, n270);
  and g313 (n271, n_224, n_225);
  not g314 (n_226, n271);
  and g315 (n272, \A[81] , n_226);
  not g316 (n_227, n268);
  not g317 (n_228, n272);
  and g318 (n273, n_227, n_228);
  not g319 (n_230, \A[79] );
  not g320 (n_231, n273);
  and g321 (n274, n_230, n_231);
  not g322 (n_233, \A[80] );
  and g323 (n275, n_233, n_226);
  and g324 (n276, \A[80] , n_231);
  not g325 (n_234, n275);
  not g326 (n_235, n276);
  and g327 (n277, n_234, n_235);
  not g328 (n_236, n277);
  and g329 (n278, \A[79] , n_236);
  not g330 (n_237, n274);
  not g331 (n_238, n278);
  and g332 (n279, n_237, n_238);
  not g333 (n_240, \A[77] );
  not g334 (n_241, n279);
  and g335 (n280, n_240, n_241);
  not g336 (n_243, \A[78] );
  and g337 (n281, n_243, n_236);
  and g338 (n282, \A[78] , n_241);
  not g339 (n_244, n281);
  not g340 (n_245, n282);
  and g341 (n283, n_244, n_245);
  not g342 (n_246, n283);
  and g343 (n284, \A[77] , n_246);
  not g344 (n_247, n280);
  not g345 (n_248, n284);
  and g346 (n285, n_247, n_248);
  not g347 (n_250, \A[75] );
  not g348 (n_251, n285);
  and g349 (n286, n_250, n_251);
  not g350 (n_253, \A[76] );
  and g351 (n287, n_253, n_246);
  and g352 (n288, \A[76] , n_251);
  not g353 (n_254, n287);
  not g354 (n_255, n288);
  and g355 (n289, n_254, n_255);
  not g356 (n_256, n289);
  and g357 (n290, \A[75] , n_256);
  not g358 (n_257, n286);
  not g359 (n_258, n290);
  and g360 (n291, n_257, n_258);
  not g361 (n_260, \A[73] );
  not g362 (n_261, n291);
  and g363 (n292, n_260, n_261);
  not g364 (n_263, \A[74] );
  and g365 (n293, n_263, n_256);
  and g366 (n294, \A[74] , n_261);
  not g367 (n_264, n293);
  not g368 (n_265, n294);
  and g369 (n295, n_264, n_265);
  not g370 (n_266, n295);
  and g371 (n296, \A[73] , n_266);
  not g372 (n_267, n292);
  not g373 (n_268, n296);
  and g374 (n297, n_267, n_268);
  not g375 (n_270, \A[71] );
  not g376 (n_271, n297);
  and g377 (n298, n_270, n_271);
  not g378 (n_273, \A[72] );
  and g379 (n299, n_273, n_266);
  and g380 (n300, \A[72] , n_271);
  not g381 (n_274, n299);
  not g382 (n_275, n300);
  and g383 (n301, n_274, n_275);
  not g384 (n_276, n301);
  and g385 (n302, \A[71] , n_276);
  not g386 (n_277, n298);
  not g387 (n_278, n302);
  and g388 (n303, n_277, n_278);
  not g389 (n_280, \A[69] );
  not g390 (n_281, n303);
  and g391 (n304, n_280, n_281);
  not g392 (n_283, \A[70] );
  and g393 (n305, n_283, n_276);
  and g394 (n306, \A[70] , n_281);
  not g395 (n_284, n305);
  not g396 (n_285, n306);
  and g397 (n307, n_284, n_285);
  not g398 (n_286, n307);
  and g399 (n308, \A[69] , n_286);
  not g400 (n_287, n304);
  not g401 (n_288, n308);
  and g402 (n309, n_287, n_288);
  not g403 (n_290, \A[67] );
  not g404 (n_291, n309);
  and g405 (n310, n_290, n_291);
  not g406 (n_293, \A[68] );
  and g407 (n311, n_293, n_286);
  and g408 (n312, \A[68] , n_291);
  not g409 (n_294, n311);
  not g410 (n_295, n312);
  and g411 (n313, n_294, n_295);
  not g412 (n_296, n313);
  and g413 (n314, \A[67] , n_296);
  not g414 (n_297, n310);
  not g415 (n_298, n314);
  and g416 (n315, n_297, n_298);
  not g417 (n_300, \A[65] );
  not g418 (n_301, n315);
  and g419 (n316, n_300, n_301);
  not g420 (n_303, \A[66] );
  and g421 (n317, n_303, n_296);
  and g422 (n318, \A[66] , n_301);
  not g423 (n_304, n317);
  not g424 (n_305, n318);
  and g425 (n319, n_304, n_305);
  not g426 (n_306, n319);
  and g427 (n320, \A[65] , n_306);
  not g428 (n_307, n316);
  not g429 (n_308, n320);
  and g430 (n321, n_307, n_308);
  not g431 (n_310, \A[63] );
  not g432 (n_311, n321);
  and g433 (n322, n_310, n_311);
  not g434 (n_313, \A[64] );
  and g435 (n323, n_313, n_306);
  and g436 (n324, \A[64] , n_311);
  not g437 (n_314, n323);
  not g438 (n_315, n324);
  and g439 (n325, n_314, n_315);
  not g440 (n_316, n325);
  and g441 (n326, \A[63] , n_316);
  not g442 (n_317, n322);
  not g443 (n_318, n326);
  and g444 (n327, n_317, n_318);
  not g445 (n_320, \A[61] );
  not g446 (n_321, n327);
  and g447 (n328, n_320, n_321);
  not g448 (n_323, \A[62] );
  and g449 (n329, n_323, n_316);
  and g450 (n330, \A[62] , n_321);
  not g451 (n_324, n329);
  not g452 (n_325, n330);
  and g453 (n331, n_324, n_325);
  not g454 (n_326, n331);
  and g455 (n332, \A[61] , n_326);
  not g456 (n_327, n328);
  not g457 (n_328, n332);
  and g458 (n333, n_327, n_328);
  not g459 (n_330, \A[59] );
  not g460 (n_331, n333);
  and g461 (n334, n_330, n_331);
  not g462 (n_333, \A[60] );
  and g463 (n335, n_333, n_326);
  and g464 (n336, \A[60] , n_331);
  not g465 (n_334, n335);
  not g466 (n_335, n336);
  and g467 (n337, n_334, n_335);
  not g468 (n_336, n337);
  and g469 (n338, \A[59] , n_336);
  not g470 (n_337, n334);
  not g471 (n_338, n338);
  and g472 (n339, n_337, n_338);
  not g473 (n_340, \A[57] );
  not g474 (n_341, n339);
  and g475 (n340, n_340, n_341);
  not g476 (n_343, \A[58] );
  and g477 (n341, n_343, n_336);
  and g478 (n342, \A[58] , n_341);
  not g479 (n_344, n341);
  not g480 (n_345, n342);
  and g481 (n343, n_344, n_345);
  not g482 (n_346, n343);
  and g483 (n344, \A[57] , n_346);
  not g484 (n_347, n340);
  not g485 (n_348, n344);
  and g486 (n345, n_347, n_348);
  not g487 (n_350, \A[55] );
  not g488 (n_351, n345);
  and g489 (n346, n_350, n_351);
  not g490 (n_353, \A[56] );
  and g491 (n347, n_353, n_346);
  and g492 (n348, \A[56] , n_351);
  not g493 (n_354, n347);
  not g494 (n_355, n348);
  and g495 (n349, n_354, n_355);
  not g496 (n_356, n349);
  and g497 (n350, \A[55] , n_356);
  not g498 (n_357, n346);
  not g499 (n_358, n350);
  and g500 (n351, n_357, n_358);
  not g501 (n_360, \A[53] );
  not g502 (n_361, n351);
  and g503 (n352, n_360, n_361);
  not g504 (n_363, \A[54] );
  and g505 (n353, n_363, n_356);
  and g506 (n354, \A[54] , n_361);
  not g507 (n_364, n353);
  not g508 (n_365, n354);
  and g509 (n355, n_364, n_365);
  not g510 (n_366, n355);
  and g511 (n356, \A[53] , n_366);
  not g512 (n_367, n352);
  not g513 (n_368, n356);
  and g514 (n357, n_367, n_368);
  not g515 (n_370, \A[51] );
  not g516 (n_371, n357);
  and g517 (n358, n_370, n_371);
  not g518 (n_373, \A[52] );
  and g519 (n359, n_373, n_366);
  and g520 (n360, \A[52] , n_371);
  not g521 (n_374, n359);
  not g522 (n_375, n360);
  and g523 (n361, n_374, n_375);
  not g524 (n_376, n361);
  and g525 (n362, \A[51] , n_376);
  not g526 (n_377, n358);
  not g527 (n_378, n362);
  and g528 (n363, n_377, n_378);
  not g529 (n_380, \A[49] );
  not g530 (n_381, n363);
  and g531 (n364, n_380, n_381);
  not g532 (n_383, \A[50] );
  and g533 (n365, n_383, n_376);
  and g534 (n366, \A[50] , n_381);
  not g535 (n_384, n365);
  not g536 (n_385, n366);
  and g537 (n367, n_384, n_385);
  not g538 (n_386, n367);
  and g539 (n368, \A[49] , n_386);
  not g540 (n_387, n364);
  not g541 (n_388, n368);
  and g542 (n369, n_387, n_388);
  not g543 (n_390, \A[47] );
  not g544 (n_391, n369);
  and g545 (n370, n_390, n_391);
  not g546 (n_393, \A[48] );
  and g547 (n371, n_393, n_386);
  and g548 (n372, \A[48] , n_391);
  not g549 (n_394, n371);
  not g550 (n_395, n372);
  and g551 (n373, n_394, n_395);
  not g552 (n_396, n373);
  and g553 (n374, \A[47] , n_396);
  not g554 (n_397, n370);
  not g555 (n_398, n374);
  and g556 (n375, n_397, n_398);
  not g557 (n_400, \A[45] );
  not g558 (n_401, n375);
  and g559 (n376, n_400, n_401);
  not g560 (n_403, \A[46] );
  and g561 (n377, n_403, n_396);
  and g562 (n378, \A[46] , n_401);
  not g563 (n_404, n377);
  not g564 (n_405, n378);
  and g565 (n379, n_404, n_405);
  not g566 (n_406, n379);
  and g567 (n380, \A[45] , n_406);
  not g568 (n_407, n376);
  not g569 (n_408, n380);
  and g570 (n381, n_407, n_408);
  not g571 (n_410, \A[43] );
  not g572 (n_411, n381);
  and g573 (n382, n_410, n_411);
  not g574 (n_413, \A[44] );
  and g575 (n383, n_413, n_406);
  and g576 (n384, \A[44] , n_411);
  not g577 (n_414, n383);
  not g578 (n_415, n384);
  and g579 (n385, n_414, n_415);
  not g580 (n_416, n385);
  and g581 (n386, \A[43] , n_416);
  not g582 (n_417, n382);
  not g583 (n_418, n386);
  and g584 (n387, n_417, n_418);
  not g585 (n_420, \A[41] );
  not g586 (n_421, n387);
  and g587 (n388, n_420, n_421);
  not g588 (n_423, \A[42] );
  and g589 (n389, n_423, n_416);
  and g590 (n390, \A[42] , n_421);
  not g591 (n_424, n389);
  not g592 (n_425, n390);
  and g593 (n391, n_424, n_425);
  not g594 (n_426, n391);
  and g595 (n392, \A[41] , n_426);
  not g596 (n_427, n388);
  not g597 (n_428, n392);
  and g598 (n393, n_427, n_428);
  not g599 (n_430, \A[39] );
  not g600 (n_431, n393);
  and g601 (n394, n_430, n_431);
  not g602 (n_433, \A[40] );
  and g603 (n395, n_433, n_426);
  and g604 (n396, \A[40] , n_431);
  not g605 (n_434, n395);
  not g606 (n_435, n396);
  and g607 (n397, n_434, n_435);
  not g608 (n_436, n397);
  and g609 (n398, \A[39] , n_436);
  not g610 (n_437, n394);
  not g611 (n_438, n398);
  and g612 (n399, n_437, n_438);
  not g613 (n_440, \A[37] );
  not g614 (n_441, n399);
  and g615 (n400, n_440, n_441);
  not g616 (n_443, \A[38] );
  and g617 (n401, n_443, n_436);
  and g618 (n402, \A[38] , n_441);
  not g619 (n_444, n401);
  not g620 (n_445, n402);
  and g621 (n403, n_444, n_445);
  not g622 (n_446, n403);
  and g623 (n404, \A[37] , n_446);
  not g624 (n_447, n400);
  not g625 (n_448, n404);
  and g626 (n405, n_447, n_448);
  not g627 (n_450, \A[35] );
  not g628 (n_451, n405);
  and g629 (n406, n_450, n_451);
  not g630 (n_453, \A[36] );
  and g631 (n407, n_453, n_446);
  and g632 (n408, \A[36] , n_451);
  not g633 (n_454, n407);
  not g634 (n_455, n408);
  and g635 (n409, n_454, n_455);
  not g636 (n_456, n409);
  and g637 (n410, \A[35] , n_456);
  not g638 (n_457, n406);
  not g639 (n_458, n410);
  and g640 (n411, n_457, n_458);
  not g641 (n_460, \A[33] );
  not g642 (n_461, n411);
  and g643 (n412, n_460, n_461);
  not g644 (n_463, \A[34] );
  and g645 (n413, n_463, n_456);
  and g646 (n414, \A[34] , n_461);
  not g647 (n_464, n413);
  not g648 (n_465, n414);
  and g649 (n415, n_464, n_465);
  not g650 (n_466, n415);
  and g651 (n416, \A[33] , n_466);
  not g652 (n_467, n412);
  not g653 (n_468, n416);
  and g654 (n417, n_467, n_468);
  not g655 (n_470, \A[31] );
  not g656 (n_471, n417);
  and g657 (n418, n_470, n_471);
  not g658 (n_473, \A[32] );
  and g659 (n419, n_473, n_466);
  and g660 (n420, \A[32] , n_471);
  not g661 (n_474, n419);
  not g662 (n_475, n420);
  and g663 (n421, n_474, n_475);
  not g664 (n_476, n421);
  and g665 (n422, \A[31] , n_476);
  not g666 (n_477, n418);
  not g667 (n_478, n422);
  and g668 (n423, n_477, n_478);
  not g669 (n_480, \A[29] );
  not g670 (n_481, n423);
  and g671 (n424, n_480, n_481);
  not g672 (n_483, \A[30] );
  and g673 (n425, n_483, n_476);
  and g674 (n426, \A[30] , n_481);
  not g675 (n_484, n425);
  not g676 (n_485, n426);
  and g677 (n427, n_484, n_485);
  not g678 (n_486, n427);
  and g679 (n428, \A[29] , n_486);
  not g680 (n_487, n424);
  not g681 (n_488, n428);
  and g682 (n429, n_487, n_488);
  not g683 (n_490, \A[27] );
  not g684 (n_491, n429);
  and g685 (n430, n_490, n_491);
  not g686 (n_493, \A[28] );
  and g687 (n431, n_493, n_486);
  and g688 (n432, \A[28] , n_491);
  not g689 (n_494, n431);
  not g690 (n_495, n432);
  and g691 (n433, n_494, n_495);
  not g692 (n_496, n433);
  and g693 (n434, \A[27] , n_496);
  not g694 (n_497, n430);
  not g695 (n_498, n434);
  and g696 (n435, n_497, n_498);
  not g697 (n_500, \A[25] );
  not g698 (n_501, n435);
  and g699 (n436, n_500, n_501);
  not g700 (n_503, \A[26] );
  and g701 (n437, n_503, n_496);
  and g702 (n438, \A[26] , n_501);
  not g703 (n_504, n437);
  not g704 (n_505, n438);
  and g705 (n439, n_504, n_505);
  not g706 (n_506, n439);
  and g707 (n440, \A[25] , n_506);
  not g708 (n_507, n436);
  not g709 (n_508, n440);
  and g710 (n441, n_507, n_508);
  not g711 (n_510, \A[23] );
  not g712 (n_511, n441);
  and g713 (n442, n_510, n_511);
  not g714 (n_513, \A[24] );
  and g715 (n443, n_513, n_506);
  and g716 (n444, \A[24] , n_511);
  not g717 (n_514, n443);
  not g718 (n_515, n444);
  and g719 (n445, n_514, n_515);
  not g720 (n_516, n445);
  and g721 (n446, \A[23] , n_516);
  not g722 (n_517, n442);
  not g723 (n_518, n446);
  and g724 (n447, n_517, n_518);
  not g725 (n_520, \A[21] );
  not g726 (n_521, n447);
  and g727 (n448, n_520, n_521);
  not g728 (n_523, \A[22] );
  and g729 (n449, n_523, n_516);
  and g730 (n450, \A[22] , n_521);
  not g731 (n_524, n449);
  not g732 (n_525, n450);
  and g733 (n451, n_524, n_525);
  not g734 (n_526, n451);
  and g735 (n452, \A[21] , n_526);
  not g736 (n_527, n448);
  not g737 (n_528, n452);
  and g738 (n453, n_527, n_528);
  not g739 (n_530, \A[19] );
  not g740 (n_531, n453);
  and g741 (n454, n_530, n_531);
  not g742 (n_533, \A[20] );
  and g743 (n455, n_533, n_526);
  and g744 (n456, \A[20] , n_531);
  not g745 (n_534, n455);
  not g746 (n_535, n456);
  and g747 (n457, n_534, n_535);
  not g748 (n_536, n457);
  and g749 (n458, \A[19] , n_536);
  not g750 (n_537, n454);
  not g751 (n_538, n458);
  and g752 (n459, n_537, n_538);
  not g753 (n_540, \A[17] );
  not g754 (n_541, n459);
  and g755 (n460, n_540, n_541);
  not g756 (n_543, \A[18] );
  and g757 (n461, n_543, n_536);
  and g758 (n462, \A[18] , n_541);
  not g759 (n_544, n461);
  not g760 (n_545, n462);
  and g761 (n463, n_544, n_545);
  not g762 (n_546, n463);
  and g763 (n464, \A[17] , n_546);
  not g764 (n_547, n460);
  not g765 (n_548, n464);
  and g766 (n465, n_547, n_548);
  not g767 (n_550, \A[15] );
  not g768 (n_551, n465);
  and g769 (n466, n_550, n_551);
  not g770 (n_553, \A[16] );
  and g771 (n467, n_553, n_546);
  and g772 (n468, \A[16] , n_551);
  not g773 (n_554, n467);
  not g774 (n_555, n468);
  and g775 (n469, n_554, n_555);
  not g776 (n_556, n469);
  and g777 (n470, \A[15] , n_556);
  not g778 (n_557, n466);
  not g779 (n_558, n470);
  and g780 (n471, n_557, n_558);
  not g781 (n_560, \A[13] );
  not g782 (n_561, n471);
  and g783 (n472, n_560, n_561);
  not g784 (n_563, \A[14] );
  and g785 (n473, n_563, n_556);
  and g786 (n474, \A[14] , n_561);
  not g787 (n_564, n473);
  not g788 (n_565, n474);
  and g789 (n475, n_564, n_565);
  not g790 (n_566, n475);
  and g791 (n476, \A[13] , n_566);
  not g792 (n_567, n472);
  not g793 (n_568, n476);
  and g794 (n477, n_567, n_568);
  not g795 (n_570, \A[11] );
  not g796 (n_571, n477);
  and g797 (n478, n_570, n_571);
  not g798 (n_573, \A[12] );
  and g799 (n479, n_573, n_566);
  and g800 (n480, \A[12] , n_571);
  not g801 (n_574, n479);
  not g802 (n_575, n480);
  and g803 (n481, n_574, n_575);
  not g804 (n_576, n481);
  and g805 (n482, \A[11] , n_576);
  not g806 (n_577, n478);
  not g807 (n_578, n482);
  and g808 (n483, n_577, n_578);
  not g809 (n_580, \A[9] );
  not g810 (n_581, n483);
  and g811 (n484, n_580, n_581);
  not g812 (n_583, \A[10] );
  and g813 (n485, n_583, n_576);
  and g814 (n486, \A[10] , n_581);
  not g815 (n_584, n485);
  not g816 (n_585, n486);
  and g817 (n487, n_584, n_585);
  not g818 (n_586, n487);
  and g819 (n488, \A[9] , n_586);
  not g820 (n_587, n484);
  not g821 (n_588, n488);
  and g822 (n489, n_587, n_588);
  not g823 (n_590, \A[7] );
  not g824 (n_591, n489);
  and g825 (n490, n_590, n_591);
  not g826 (n_593, \A[8] );
  and g827 (n491, n_593, n_586);
  and g828 (n492, \A[8] , n_591);
  not g829 (n_594, n491);
  not g830 (n_595, n492);
  and g831 (n493, n_594, n_595);
  not g832 (n_596, n493);
  and g833 (n494, \A[7] , n_596);
  not g834 (n_597, n490);
  not g835 (n_598, n494);
  and g836 (n495, n_597, n_598);
  not g837 (n_600, \A[5] );
  not g838 (n_601, n495);
  and g839 (n496, n_600, n_601);
  not g840 (n_603, \A[6] );
  and g841 (n497, n_603, n_596);
  and g842 (n498, \A[6] , n_601);
  not g843 (n_604, n497);
  not g844 (n_605, n498);
  and g845 (n499, n_604, n_605);
  not g846 (n_606, n499);
  and g847 (n500, \A[5] , n_606);
  not g848 (n_607, n496);
  not g849 (n_608, n500);
  and g850 (n501, n_607, n_608);
  not g851 (n_610, \A[3] );
  not g852 (n_611, n501);
  and g853 (n502, n_610, n_611);
  not g854 (n_613, \A[4] );
  and g855 (n503, n_613, n_606);
  and g856 (n504, \A[4] , n_611);
  not g857 (n_614, n503);
  not g858 (n_615, n504);
  and g859 (n505, n_614, n_615);
  not g860 (n_616, n505);
  and g861 (n506, \A[3] , n_616);
  not g862 (n_617, n502);
  not g863 (n_618, n506);
  and g864 (n507, n_617, n_618);
  not g865 (n_621, \A[2] );
  and g866 (n508, \A[1] , n_621);
  not g867 (n_622, n508);
  and g868 (n509, n507, n_622);
  and g869 (n510, n505, n508);
  not g870 (n_623, n509);
  not g871 (n_624, n510);
  and g872 (\P[0] , n_623, n_624);
  not g873 (n_625, \A[126] );
  and g874 (n512, n_625, \A[127] );
  not g875 (n_626, n512);
  and g876 (n513, n_625, n_626);
  and g877 (n514, n_13, n_2);
  and g878 (n515, n_23, n_10);
  and g879 (n516, \A[121] , n515);
  not g880 (n_627, n516);
  and g881 (n517, n514, n_627);
  not g882 (n_628, n517);
  and g883 (n518, n513, n_628);
  not g884 (n_629, n518);
  and g885 (n519, n_33, n_629);
  not g886 (n_630, n515);
  and g887 (n520, n514, n_630);
  not g888 (n_631, n520);
  and g889 (n521, n513, n_631);
  not g890 (n_632, n521);
  and g891 (n522, \A[120] , n_632);
  not g892 (n_633, n519);
  not g893 (n_634, n522);
  and g894 (n523, n_633, n_634);
  and g895 (n524, n_43, n_30);
  not g896 (n_635, n524);
  and g897 (n525, n523, n_635);
  and g898 (n526, n521, n524);
  not g899 (n_636, n525);
  not g900 (n_637, n526);
  and g901 (n527, n_636, n_637);
  and g902 (n528, n_53, n_40);
  not g903 (n_638, n528);
  and g904 (n529, n527, n_638);
  not g905 (n_639, n523);
  and g906 (n530, n_639, n528);
  not g907 (n_640, n529);
  not g908 (n_641, n530);
  and g909 (n531, n_640, n_641);
  and g910 (n532, n_63, n_50);
  not g911 (n_642, n532);
  and g912 (n533, n531, n_642);
  not g913 (n_643, n527);
  and g914 (n534, n_643, n532);
  not g915 (n_644, n533);
  not g916 (n_645, n534);
  and g917 (n535, n_644, n_645);
  and g918 (n536, n_73, n_60);
  not g919 (n_646, n536);
  and g920 (n537, n535, n_646);
  not g921 (n_647, n531);
  and g922 (n538, n_647, n536);
  not g923 (n_648, n537);
  not g924 (n_649, n538);
  and g925 (n539, n_648, n_649);
  and g926 (n540, n_83, n_70);
  not g927 (n_650, n540);
  and g928 (n541, n539, n_650);
  not g929 (n_651, n535);
  and g930 (n542, n_651, n540);
  not g931 (n_652, n541);
  not g932 (n_653, n542);
  and g933 (n543, n_652, n_653);
  and g934 (n544, n_93, n_80);
  not g935 (n_654, n544);
  and g936 (n545, n543, n_654);
  not g937 (n_655, n539);
  and g938 (n546, n_655, n544);
  not g939 (n_656, n545);
  not g940 (n_657, n546);
  and g941 (n547, n_656, n_657);
  and g942 (n548, n_103, n_90);
  not g943 (n_658, n548);
  and g944 (n549, n547, n_658);
  not g945 (n_659, n543);
  and g946 (n550, n_659, n548);
  not g947 (n_660, n549);
  not g948 (n_661, n550);
  and g949 (n551, n_660, n_661);
  and g950 (n552, n_113, n_100);
  not g951 (n_662, n552);
  and g952 (n553, n551, n_662);
  not g953 (n_663, n547);
  and g954 (n554, n_663, n552);
  not g955 (n_664, n553);
  not g956 (n_665, n554);
  and g957 (n555, n_664, n_665);
  and g958 (n556, n_123, n_110);
  not g959 (n_666, n556);
  and g960 (n557, n555, n_666);
  not g961 (n_667, n551);
  and g962 (n558, n_667, n556);
  not g963 (n_668, n557);
  not g964 (n_669, n558);
  and g965 (n559, n_668, n_669);
  and g966 (n560, n_133, n_120);
  not g967 (n_670, n560);
  and g968 (n561, n559, n_670);
  not g969 (n_671, n555);
  and g970 (n562, n_671, n560);
  not g971 (n_672, n561);
  not g972 (n_673, n562);
  and g973 (n563, n_672, n_673);
  and g974 (n564, n_143, n_130);
  not g975 (n_674, n564);
  and g976 (n565, n563, n_674);
  not g977 (n_675, n559);
  and g978 (n566, n_675, n564);
  not g979 (n_676, n565);
  not g980 (n_677, n566);
  and g981 (n567, n_676, n_677);
  and g982 (n568, n_153, n_140);
  not g983 (n_678, n568);
  and g984 (n569, n567, n_678);
  not g985 (n_679, n563);
  and g986 (n570, n_679, n568);
  not g987 (n_680, n569);
  not g988 (n_681, n570);
  and g989 (n571, n_680, n_681);
  and g990 (n572, n_163, n_150);
  not g991 (n_682, n572);
  and g992 (n573, n571, n_682);
  not g993 (n_683, n567);
  and g994 (n574, n_683, n572);
  not g995 (n_684, n573);
  not g996 (n_685, n574);
  and g997 (n575, n_684, n_685);
  and g998 (n576, n_173, n_160);
  not g999 (n_686, n576);
  and g1000 (n577, n575, n_686);
  not g1001 (n_687, n571);
  and g1002 (n578, n_687, n576);
  not g1003 (n_688, n577);
  not g1004 (n_689, n578);
  and g1005 (n579, n_688, n_689);
  and g1006 (n580, n_183, n_170);
  not g1007 (n_690, n580);
  and g1008 (n581, n579, n_690);
  not g1009 (n_691, n575);
  and g1010 (n582, n_691, n580);
  not g1011 (n_692, n581);
  not g1012 (n_693, n582);
  and g1013 (n583, n_692, n_693);
  and g1014 (n584, n_193, n_180);
  not g1015 (n_694, n584);
  and g1016 (n585, n583, n_694);
  not g1017 (n_695, n579);
  and g1018 (n586, n_695, n584);
  not g1019 (n_696, n585);
  not g1020 (n_697, n586);
  and g1021 (n587, n_696, n_697);
  and g1022 (n588, n_203, n_190);
  not g1023 (n_698, n588);
  and g1024 (n589, n587, n_698);
  not g1025 (n_699, n583);
  and g1026 (n590, n_699, n588);
  not g1027 (n_700, n589);
  not g1028 (n_701, n590);
  and g1029 (n591, n_700, n_701);
  and g1030 (n592, n_213, n_200);
  not g1031 (n_702, n592);
  and g1032 (n593, n591, n_702);
  not g1033 (n_703, n587);
  and g1034 (n594, n_703, n592);
  not g1035 (n_704, n593);
  not g1036 (n_705, n594);
  and g1037 (n595, n_704, n_705);
  and g1038 (n596, n_223, n_210);
  not g1039 (n_706, n596);
  and g1040 (n597, n595, n_706);
  not g1041 (n_707, n591);
  and g1042 (n598, n_707, n596);
  not g1043 (n_708, n597);
  not g1044 (n_709, n598);
  and g1045 (n599, n_708, n_709);
  and g1046 (n600, n_233, n_220);
  not g1047 (n_710, n600);
  and g1048 (n601, n599, n_710);
  not g1049 (n_711, n595);
  and g1050 (n602, n_711, n600);
  not g1051 (n_712, n601);
  not g1052 (n_713, n602);
  and g1053 (n603, n_712, n_713);
  and g1054 (n604, n_243, n_230);
  not g1055 (n_714, n604);
  and g1056 (n605, n603, n_714);
  not g1057 (n_715, n599);
  and g1058 (n606, n_715, n604);
  not g1059 (n_716, n605);
  not g1060 (n_717, n606);
  and g1061 (n607, n_716, n_717);
  and g1062 (n608, n_253, n_240);
  not g1063 (n_718, n608);
  and g1064 (n609, n607, n_718);
  not g1065 (n_719, n603);
  and g1066 (n610, n_719, n608);
  not g1067 (n_720, n609);
  not g1068 (n_721, n610);
  and g1069 (n611, n_720, n_721);
  and g1070 (n612, n_263, n_250);
  not g1071 (n_722, n612);
  and g1072 (n613, n611, n_722);
  not g1073 (n_723, n607);
  and g1074 (n614, n_723, n612);
  not g1075 (n_724, n613);
  not g1076 (n_725, n614);
  and g1077 (n615, n_724, n_725);
  and g1078 (n616, n_273, n_260);
  not g1079 (n_726, n616);
  and g1080 (n617, n615, n_726);
  not g1081 (n_727, n611);
  and g1082 (n618, n_727, n616);
  not g1083 (n_728, n617);
  not g1084 (n_729, n618);
  and g1085 (n619, n_728, n_729);
  and g1086 (n620, n_283, n_270);
  not g1087 (n_730, n620);
  and g1088 (n621, n619, n_730);
  not g1089 (n_731, n615);
  and g1090 (n622, n_731, n620);
  not g1091 (n_732, n621);
  not g1092 (n_733, n622);
  and g1093 (n623, n_732, n_733);
  and g1094 (n624, n_293, n_280);
  not g1095 (n_734, n624);
  and g1096 (n625, n623, n_734);
  not g1097 (n_735, n619);
  and g1098 (n626, n_735, n624);
  not g1099 (n_736, n625);
  not g1100 (n_737, n626);
  and g1101 (n627, n_736, n_737);
  and g1102 (n628, n_303, n_290);
  not g1103 (n_738, n628);
  and g1104 (n629, n627, n_738);
  not g1105 (n_739, n623);
  and g1106 (n630, n_739, n628);
  not g1107 (n_740, n629);
  not g1108 (n_741, n630);
  and g1109 (n631, n_740, n_741);
  and g1110 (n632, n_313, n_300);
  not g1111 (n_742, n632);
  and g1112 (n633, n631, n_742);
  not g1113 (n_743, n627);
  and g1114 (n634, n_743, n632);
  not g1115 (n_744, n633);
  not g1116 (n_745, n634);
  and g1117 (n635, n_744, n_745);
  and g1118 (n636, n_323, n_310);
  not g1119 (n_746, n636);
  and g1120 (n637, n635, n_746);
  not g1121 (n_747, n631);
  and g1122 (n638, n_747, n636);
  not g1123 (n_748, n637);
  not g1124 (n_749, n638);
  and g1125 (n639, n_748, n_749);
  and g1126 (n640, n_333, n_320);
  not g1127 (n_750, n640);
  and g1128 (n641, n639, n_750);
  not g1129 (n_751, n635);
  and g1130 (n642, n_751, n640);
  not g1131 (n_752, n641);
  not g1132 (n_753, n642);
  and g1133 (n643, n_752, n_753);
  and g1134 (n644, n_343, n_330);
  not g1135 (n_754, n644);
  and g1136 (n645, n643, n_754);
  not g1137 (n_755, n639);
  and g1138 (n646, n_755, n644);
  not g1139 (n_756, n645);
  not g1140 (n_757, n646);
  and g1141 (n647, n_756, n_757);
  and g1142 (n648, n_353, n_340);
  not g1143 (n_758, n648);
  and g1144 (n649, n647, n_758);
  not g1145 (n_759, n643);
  and g1146 (n650, n_759, n648);
  not g1147 (n_760, n649);
  not g1148 (n_761, n650);
  and g1149 (n651, n_760, n_761);
  and g1150 (n652, n_363, n_350);
  not g1151 (n_762, n652);
  and g1152 (n653, n651, n_762);
  not g1153 (n_763, n647);
  and g1154 (n654, n_763, n652);
  not g1155 (n_764, n653);
  not g1156 (n_765, n654);
  and g1157 (n655, n_764, n_765);
  and g1158 (n656, n_373, n_360);
  not g1159 (n_766, n656);
  and g1160 (n657, n655, n_766);
  not g1161 (n_767, n651);
  and g1162 (n658, n_767, n656);
  not g1163 (n_768, n657);
  not g1164 (n_769, n658);
  and g1165 (n659, n_768, n_769);
  and g1166 (n660, n_383, n_370);
  not g1167 (n_770, n660);
  and g1168 (n661, n659, n_770);
  not g1169 (n_771, n655);
  and g1170 (n662, n_771, n660);
  not g1171 (n_772, n661);
  not g1172 (n_773, n662);
  and g1173 (n663, n_772, n_773);
  and g1174 (n664, n_393, n_380);
  not g1175 (n_774, n664);
  and g1176 (n665, n663, n_774);
  not g1177 (n_775, n659);
  and g1178 (n666, n_775, n664);
  not g1179 (n_776, n665);
  not g1180 (n_777, n666);
  and g1181 (n667, n_776, n_777);
  and g1182 (n668, n_403, n_390);
  not g1183 (n_778, n668);
  and g1184 (n669, n667, n_778);
  not g1185 (n_779, n663);
  and g1186 (n670, n_779, n668);
  not g1187 (n_780, n669);
  not g1188 (n_781, n670);
  and g1189 (n671, n_780, n_781);
  and g1190 (n672, n_413, n_400);
  not g1191 (n_782, n672);
  and g1192 (n673, n671, n_782);
  not g1193 (n_783, n667);
  and g1194 (n674, n_783, n672);
  not g1195 (n_784, n673);
  not g1196 (n_785, n674);
  and g1197 (n675, n_784, n_785);
  and g1198 (n676, n_423, n_410);
  not g1199 (n_786, n676);
  and g1200 (n677, n675, n_786);
  not g1201 (n_787, n671);
  and g1202 (n678, n_787, n676);
  not g1203 (n_788, n677);
  not g1204 (n_789, n678);
  and g1205 (n679, n_788, n_789);
  and g1206 (n680, n_433, n_420);
  not g1207 (n_790, n680);
  and g1208 (n681, n679, n_790);
  not g1209 (n_791, n675);
  and g1210 (n682, n_791, n680);
  not g1211 (n_792, n681);
  not g1212 (n_793, n682);
  and g1213 (n683, n_792, n_793);
  and g1214 (n684, n_443, n_430);
  not g1215 (n_794, n684);
  and g1216 (n685, n683, n_794);
  not g1217 (n_795, n679);
  and g1218 (n686, n_795, n684);
  not g1219 (n_796, n685);
  not g1220 (n_797, n686);
  and g1221 (n687, n_796, n_797);
  and g1222 (n688, n_453, n_440);
  not g1223 (n_798, n688);
  and g1224 (n689, n687, n_798);
  not g1225 (n_799, n683);
  and g1226 (n690, n_799, n688);
  not g1227 (n_800, n689);
  not g1228 (n_801, n690);
  and g1229 (n691, n_800, n_801);
  and g1230 (n692, n_463, n_450);
  not g1231 (n_802, n692);
  and g1232 (n693, n691, n_802);
  not g1233 (n_803, n687);
  and g1234 (n694, n_803, n692);
  not g1235 (n_804, n693);
  not g1236 (n_805, n694);
  and g1237 (n695, n_804, n_805);
  and g1238 (n696, n_473, n_460);
  not g1239 (n_806, n696);
  and g1240 (n697, n695, n_806);
  not g1241 (n_807, n691);
  and g1242 (n698, n_807, n696);
  not g1243 (n_808, n697);
  not g1244 (n_809, n698);
  and g1245 (n699, n_808, n_809);
  and g1246 (n700, n_483, n_470);
  not g1247 (n_810, n700);
  and g1248 (n701, n699, n_810);
  not g1249 (n_811, n695);
  and g1250 (n702, n_811, n700);
  not g1251 (n_812, n701);
  not g1252 (n_813, n702);
  and g1253 (n703, n_812, n_813);
  and g1254 (n704, n_493, n_480);
  not g1255 (n_814, n704);
  and g1256 (n705, n703, n_814);
  not g1257 (n_815, n699);
  and g1258 (n706, n_815, n704);
  not g1259 (n_816, n705);
  not g1260 (n_817, n706);
  and g1261 (n707, n_816, n_817);
  and g1262 (n708, n_503, n_490);
  not g1263 (n_818, n708);
  and g1264 (n709, n707, n_818);
  not g1265 (n_819, n703);
  and g1266 (n710, n_819, n708);
  not g1267 (n_820, n709);
  not g1268 (n_821, n710);
  and g1269 (n711, n_820, n_821);
  and g1270 (n712, n_513, n_500);
  not g1271 (n_822, n712);
  and g1272 (n713, n711, n_822);
  not g1273 (n_823, n707);
  and g1274 (n714, n_823, n712);
  not g1275 (n_824, n713);
  not g1276 (n_825, n714);
  and g1277 (n715, n_824, n_825);
  and g1278 (n716, n_523, n_510);
  not g1279 (n_826, n716);
  and g1280 (n717, n715, n_826);
  not g1281 (n_827, n711);
  and g1282 (n718, n_827, n716);
  not g1283 (n_828, n717);
  not g1284 (n_829, n718);
  and g1285 (n719, n_828, n_829);
  and g1286 (n720, n_533, n_520);
  not g1287 (n_830, n720);
  and g1288 (n721, n719, n_830);
  not g1289 (n_831, n715);
  and g1290 (n722, n_831, n720);
  not g1291 (n_832, n721);
  not g1292 (n_833, n722);
  and g1293 (n723, n_832, n_833);
  and g1294 (n724, n_543, n_530);
  not g1295 (n_834, n724);
  and g1296 (n725, n723, n_834);
  not g1297 (n_835, n719);
  and g1298 (n726, n_835, n724);
  not g1299 (n_836, n725);
  not g1300 (n_837, n726);
  and g1301 (n727, n_836, n_837);
  and g1302 (n728, n_553, n_540);
  not g1303 (n_838, n728);
  and g1304 (n729, n727, n_838);
  not g1305 (n_839, n723);
  and g1306 (n730, n_839, n728);
  not g1307 (n_840, n729);
  not g1308 (n_841, n730);
  and g1309 (n731, n_840, n_841);
  and g1310 (n732, n_563, n_550);
  not g1311 (n_842, n732);
  and g1312 (n733, n731, n_842);
  not g1313 (n_843, n727);
  and g1314 (n734, n_843, n732);
  not g1315 (n_844, n733);
  not g1316 (n_845, n734);
  and g1317 (n735, n_844, n_845);
  and g1318 (n736, n_573, n_560);
  not g1319 (n_846, n736);
  and g1320 (n737, n735, n_846);
  not g1321 (n_847, n731);
  and g1322 (n738, n_847, n736);
  not g1323 (n_848, n737);
  not g1324 (n_849, n738);
  and g1325 (n739, n_848, n_849);
  and g1326 (n740, n_583, n_570);
  not g1327 (n_850, n740);
  and g1328 (n741, n739, n_850);
  not g1329 (n_851, n735);
  and g1330 (n742, n_851, n740);
  not g1331 (n_852, n741);
  not g1332 (n_853, n742);
  and g1333 (n743, n_852, n_853);
  and g1334 (n744, n_593, n_580);
  not g1335 (n_854, n744);
  and g1336 (n745, n743, n_854);
  not g1337 (n_855, n739);
  and g1338 (n746, n_855, n744);
  not g1339 (n_856, n745);
  not g1340 (n_857, n746);
  and g1341 (n747, n_856, n_857);
  and g1342 (n748, n_603, n_590);
  not g1343 (n_858, n748);
  and g1344 (n749, n747, n_858);
  not g1345 (n_859, n743);
  and g1346 (n750, n_859, n748);
  not g1347 (n_860, n749);
  not g1348 (n_861, n750);
  and g1349 (n751, n_860, n_861);
  and g1350 (n752, n_613, n_600);
  not g1351 (n_862, n752);
  and g1352 (n753, n751, n_862);
  not g1353 (n_863, n747);
  and g1354 (n754, n_863, n752);
  not g1355 (n_864, n753);
  not g1356 (n_865, n754);
  and g1357 (n755, n_864, n_865);
  and g1358 (n756, n_621, n_610);
  not g1359 (n_866, n756);
  and g1360 (n757, n755, n_866);
  not g1361 (n_867, n751);
  and g1362 (n758, n_867, n756);
  not g1363 (n_868, n757);
  not g1364 (n_869, n758);
  and g1365 (\P[1] , n_868, n_869);
  and g1366 (n760, n513, n514);
  and g1367 (n761, n_33, n_20);
  and g1368 (n762, n515, n761);
  and g1369 (n763, n_40, n524);
  and g1370 (n764, n_53, n763);
  not g1371 (n_870, n764);
  and g1372 (n765, n762, n_870);
  not g1373 (n_871, n765);
  and g1374 (n766, n760, n_871);
  and g1375 (n767, n_60, n_63);
  and g1376 (n768, n_73, n767);
  not g1377 (n_872, n768);
  and g1378 (n769, n766, n_872);
  and g1379 (n770, \A[115] , n764);
  not g1380 (n_873, n770);
  and g1381 (n771, n762, n_873);
  not g1382 (n_874, n771);
  and g1383 (n772, n760, n_874);
  and g1384 (n773, n768, n772);
  not g1385 (n_875, n769);
  not g1386 (n_876, n773);
  and g1387 (n774, n_875, n_876);
  and g1388 (n775, n_80, n540);
  and g1389 (n776, n_93, n775);
  not g1390 (n_877, n776);
  and g1391 (n777, n774, n_877);
  not g1392 (n_878, n766);
  and g1393 (n778, n_878, n776);
  not g1394 (n_879, n777);
  not g1395 (n_880, n778);
  and g1396 (n779, n_879, n_880);
  and g1397 (n780, n_100, n548);
  and g1398 (n781, n_113, n780);
  not g1399 (n_881, n781);
  and g1400 (n782, n779, n_881);
  not g1401 (n_882, n774);
  and g1402 (n783, n_882, n781);
  not g1403 (n_883, n782);
  not g1404 (n_884, n783);
  and g1405 (n784, n_883, n_884);
  and g1406 (n785, n_120, n556);
  and g1407 (n786, n_133, n785);
  not g1408 (n_885, n786);
  and g1409 (n787, n784, n_885);
  not g1410 (n_886, n779);
  and g1411 (n788, n_886, n786);
  not g1412 (n_887, n787);
  not g1413 (n_888, n788);
  and g1414 (n789, n_887, n_888);
  and g1415 (n790, n_140, n564);
  and g1416 (n791, n_153, n790);
  not g1417 (n_889, n791);
  and g1418 (n792, n789, n_889);
  not g1419 (n_890, n784);
  and g1420 (n793, n_890, n791);
  not g1421 (n_891, n792);
  not g1422 (n_892, n793);
  and g1423 (n794, n_891, n_892);
  and g1424 (n795, n_160, n572);
  and g1425 (n796, n_173, n795);
  not g1426 (n_893, n796);
  and g1427 (n797, n794, n_893);
  not g1428 (n_894, n789);
  and g1429 (n798, n_894, n796);
  not g1430 (n_895, n797);
  not g1431 (n_896, n798);
  and g1432 (n799, n_895, n_896);
  and g1433 (n800, n_180, n580);
  and g1434 (n801, n_193, n800);
  not g1435 (n_897, n801);
  and g1436 (n802, n799, n_897);
  not g1437 (n_898, n794);
  and g1438 (n803, n_898, n801);
  not g1439 (n_899, n802);
  not g1440 (n_900, n803);
  and g1441 (n804, n_899, n_900);
  and g1442 (n805, n_200, n588);
  and g1443 (n806, n_213, n805);
  not g1444 (n_901, n806);
  and g1445 (n807, n804, n_901);
  not g1446 (n_902, n799);
  and g1447 (n808, n_902, n806);
  not g1448 (n_903, n807);
  not g1449 (n_904, n808);
  and g1450 (n809, n_903, n_904);
  and g1451 (n810, n_220, n596);
  and g1452 (n811, n_233, n810);
  not g1453 (n_905, n811);
  and g1454 (n812, n809, n_905);
  not g1455 (n_906, n804);
  and g1456 (n813, n_906, n811);
  not g1457 (n_907, n812);
  not g1458 (n_908, n813);
  and g1459 (n814, n_907, n_908);
  and g1460 (n815, n_240, n604);
  and g1461 (n816, n_253, n815);
  not g1462 (n_909, n816);
  and g1463 (n817, n814, n_909);
  not g1464 (n_910, n809);
  and g1465 (n818, n_910, n816);
  not g1466 (n_911, n817);
  not g1467 (n_912, n818);
  and g1468 (n819, n_911, n_912);
  and g1469 (n820, n_260, n612);
  and g1470 (n821, n_273, n820);
  not g1471 (n_913, n821);
  and g1472 (n822, n819, n_913);
  not g1473 (n_914, n814);
  and g1474 (n823, n_914, n821);
  not g1475 (n_915, n822);
  not g1476 (n_916, n823);
  and g1477 (n824, n_915, n_916);
  and g1478 (n825, n_280, n620);
  and g1479 (n826, n_293, n825);
  not g1480 (n_917, n826);
  and g1481 (n827, n824, n_917);
  not g1482 (n_918, n819);
  and g1483 (n828, n_918, n826);
  not g1484 (n_919, n827);
  not g1485 (n_920, n828);
  and g1486 (n829, n_919, n_920);
  and g1487 (n830, n_300, n628);
  and g1488 (n831, n_313, n830);
  not g1489 (n_921, n831);
  and g1490 (n832, n829, n_921);
  not g1491 (n_922, n824);
  and g1492 (n833, n_922, n831);
  not g1493 (n_923, n832);
  not g1494 (n_924, n833);
  and g1495 (n834, n_923, n_924);
  and g1496 (n835, n_320, n636);
  and g1497 (n836, n_333, n835);
  not g1498 (n_925, n836);
  and g1499 (n837, n834, n_925);
  not g1500 (n_926, n829);
  and g1501 (n838, n_926, n836);
  not g1502 (n_927, n837);
  not g1503 (n_928, n838);
  and g1504 (n839, n_927, n_928);
  and g1505 (n840, n_340, n644);
  and g1506 (n841, n_353, n840);
  not g1507 (n_929, n841);
  and g1508 (n842, n839, n_929);
  not g1509 (n_930, n834);
  and g1510 (n843, n_930, n841);
  not g1511 (n_931, n842);
  not g1512 (n_932, n843);
  and g1513 (n844, n_931, n_932);
  and g1514 (n845, n_360, n652);
  and g1515 (n846, n_373, n845);
  not g1516 (n_933, n846);
  and g1517 (n847, n844, n_933);
  not g1518 (n_934, n839);
  and g1519 (n848, n_934, n846);
  not g1520 (n_935, n847);
  not g1521 (n_936, n848);
  and g1522 (n849, n_935, n_936);
  and g1523 (n850, n_380, n660);
  and g1524 (n851, n_393, n850);
  not g1525 (n_937, n851);
  and g1526 (n852, n849, n_937);
  not g1527 (n_938, n844);
  and g1528 (n853, n_938, n851);
  not g1529 (n_939, n852);
  not g1530 (n_940, n853);
  and g1531 (n854, n_939, n_940);
  and g1532 (n855, n_400, n668);
  and g1533 (n856, n_413, n855);
  not g1534 (n_941, n856);
  and g1535 (n857, n854, n_941);
  not g1536 (n_942, n849);
  and g1537 (n858, n_942, n856);
  not g1538 (n_943, n857);
  not g1539 (n_944, n858);
  and g1540 (n859, n_943, n_944);
  and g1541 (n860, n_420, n676);
  and g1542 (n861, n_433, n860);
  not g1543 (n_945, n861);
  and g1544 (n862, n859, n_945);
  not g1545 (n_946, n854);
  and g1546 (n863, n_946, n861);
  not g1547 (n_947, n862);
  not g1548 (n_948, n863);
  and g1549 (n864, n_947, n_948);
  and g1550 (n865, n_440, n684);
  and g1551 (n866, n_453, n865);
  not g1552 (n_949, n866);
  and g1553 (n867, n864, n_949);
  not g1554 (n_950, n859);
  and g1555 (n868, n_950, n866);
  not g1556 (n_951, n867);
  not g1557 (n_952, n868);
  and g1558 (n869, n_951, n_952);
  and g1559 (n870, n_460, n692);
  and g1560 (n871, n_473, n870);
  not g1561 (n_953, n871);
  and g1562 (n872, n869, n_953);
  not g1563 (n_954, n864);
  and g1564 (n873, n_954, n871);
  not g1565 (n_955, n872);
  not g1566 (n_956, n873);
  and g1567 (n874, n_955, n_956);
  and g1568 (n875, n_480, n700);
  and g1569 (n876, n_493, n875);
  not g1570 (n_957, n876);
  and g1571 (n877, n874, n_957);
  not g1572 (n_958, n869);
  and g1573 (n878, n_958, n876);
  not g1574 (n_959, n877);
  not g1575 (n_960, n878);
  and g1576 (n879, n_959, n_960);
  and g1577 (n880, n_500, n708);
  and g1578 (n881, n_513, n880);
  not g1579 (n_961, n881);
  and g1580 (n882, n879, n_961);
  not g1581 (n_962, n874);
  and g1582 (n883, n_962, n881);
  not g1583 (n_963, n882);
  not g1584 (n_964, n883);
  and g1585 (n884, n_963, n_964);
  and g1586 (n885, n_520, n716);
  and g1587 (n886, n_533, n885);
  not g1588 (n_965, n886);
  and g1589 (n887, n884, n_965);
  not g1590 (n_966, n879);
  and g1591 (n888, n_966, n886);
  not g1592 (n_967, n887);
  not g1593 (n_968, n888);
  and g1594 (n889, n_967, n_968);
  and g1595 (n890, n_540, n724);
  and g1596 (n891, n_553, n890);
  not g1597 (n_969, n891);
  and g1598 (n892, n889, n_969);
  not g1599 (n_970, n884);
  and g1600 (n893, n_970, n891);
  not g1601 (n_971, n892);
  not g1602 (n_972, n893);
  and g1603 (n894, n_971, n_972);
  and g1604 (n895, n_560, n732);
  and g1605 (n896, n_573, n895);
  not g1606 (n_973, n896);
  and g1607 (n897, n894, n_973);
  not g1608 (n_974, n889);
  and g1609 (n898, n_974, n896);
  not g1610 (n_975, n897);
  not g1611 (n_976, n898);
  and g1612 (n899, n_975, n_976);
  and g1613 (n900, n_580, n740);
  and g1614 (n901, n_593, n900);
  not g1615 (n_977, n901);
  and g1616 (n902, n899, n_977);
  not g1617 (n_978, n894);
  and g1618 (n903, n_978, n901);
  not g1619 (n_979, n902);
  not g1620 (n_980, n903);
  and g1621 (n904, n_979, n_980);
  and g1622 (n905, n_600, n748);
  and g1623 (n906, n_613, n905);
  not g1624 (n_981, n906);
  and g1625 (n907, n904, n_981);
  not g1626 (n_982, n899);
  and g1627 (n908, n_982, n906);
  or g1628 (\P[2] , n907, n908);
  and g1629 (n910, n760, n762);
  not g1637 (n_983, n917);
  and g1638 (n918, n913, n_983);
  not g1639 (n_984, n918);
  and g1640 (n919, n910, n_984);
  not g1647 (n_985, n925);
  and g1648 (n926, n919, n_985);
  and g1649 (n927, \A[103] , n917);
  not g1650 (n_986, n927);
  and g1651 (n928, n913, n_986);
  not g1652 (n_987, n928);
  and g1653 (n929, n910, n_987);
  and g1654 (n930, n925, n929);
  not g1655 (n_988, n926);
  not g1656 (n_989, n930);
  and g1657 (n931, n_988, n_989);
  not g1662 (n_990, n935);
  and g1663 (n936, n931, n_990);
  not g1664 (n_991, n919);
  and g1665 (n937, n_991, n935);
  not g1666 (n_992, n936);
  not g1667 (n_993, n937);
  and g1668 (n938, n_992, n_993);
  not g1673 (n_994, n942);
  and g1674 (n943, n938, n_994);
  not g1675 (n_995, n931);
  and g1676 (n944, n_995, n942);
  not g1677 (n_996, n943);
  not g1678 (n_997, n944);
  and g1679 (n945, n_996, n_997);
  not g1684 (n_998, n949);
  and g1685 (n950, n945, n_998);
  not g1686 (n_999, n938);
  and g1687 (n951, n_999, n949);
  not g1688 (n_1000, n950);
  not g1689 (n_1001, n951);
  and g1690 (n952, n_1000, n_1001);
  not g1695 (n_1002, n956);
  and g1696 (n957, n952, n_1002);
  not g1697 (n_1003, n945);
  and g1698 (n958, n_1003, n956);
  not g1699 (n_1004, n957);
  not g1700 (n_1005, n958);
  and g1701 (n959, n_1004, n_1005);
  not g1706 (n_1006, n963);
  and g1707 (n964, n959, n_1006);
  not g1708 (n_1007, n952);
  and g1709 (n965, n_1007, n963);
  not g1710 (n_1008, n964);
  not g1711 (n_1009, n965);
  and g1712 (n966, n_1008, n_1009);
  not g1717 (n_1010, n970);
  and g1718 (n971, n966, n_1010);
  not g1719 (n_1011, n959);
  and g1720 (n972, n_1011, n970);
  not g1721 (n_1012, n971);
  not g1722 (n_1013, n972);
  and g1723 (n973, n_1012, n_1013);
  not g1728 (n_1014, n977);
  and g1729 (n978, n973, n_1014);
  not g1730 (n_1015, n966);
  and g1731 (n979, n_1015, n977);
  not g1732 (n_1016, n978);
  not g1733 (n_1017, n979);
  and g1734 (n980, n_1016, n_1017);
  not g1739 (n_1018, n984);
  and g1740 (n985, n980, n_1018);
  not g1741 (n_1019, n973);
  and g1742 (n986, n_1019, n984);
  not g1743 (n_1020, n985);
  not g1744 (n_1021, n986);
  and g1745 (n987, n_1020, n_1021);
  not g1750 (n_1022, n991);
  and g1751 (n992, n987, n_1022);
  not g1752 (n_1023, n980);
  and g1753 (n993, n_1023, n991);
  not g1754 (n_1024, n992);
  not g1755 (n_1025, n993);
  and g1756 (n994, n_1024, n_1025);
  not g1761 (n_1026, n998);
  and g1762 (n999, n994, n_1026);
  not g1763 (n_1027, n987);
  and g1764 (n1000, n_1027, n998);
  not g1765 (n_1028, n999);
  not g1766 (n_1029, n1000);
  and g1767 (n1001, n_1028, n_1029);
  not g1772 (n_1030, n1005);
  and g1773 (n1006, n1001, n_1030);
  not g1774 (n_1031, n994);
  and g1775 (n1007, n_1031, n1005);
  or g1776 (\P[3] , n1006, n1007);
  and g1777 (n1009, n910, n913);
  not g1791 (n_1032, n1022);
  and g1792 (n1023, n1014, n_1032);
  not g1793 (n_1033, n1023);
  and g1794 (n1024, n1009, n_1033);
  not g1809 (n_1034, n1038);
  and g1810 (n1039, n1024, n_1034);
  and g1811 (n1040, \A[79] , n1022);
  not g1812 (n_1035, n1040);
  and g1813 (n1041, n1014, n_1035);
  not g1814 (n_1036, n1041);
  and g1815 (n1042, n1009, n_1036);
  and g1816 (n1043, n1038, n1042);
  not g1817 (n_1037, n1039);
  not g1818 (n_1038, n1043);
  and g1819 (n1044, n_1037, n_1038);
  not g1828 (n_1039, n1052);
  and g1829 (n1053, n1044, n_1039);
  not g1830 (n_1040, n1024);
  and g1831 (n1054, n_1040, n1052);
  not g1832 (n_1041, n1053);
  not g1833 (n_1042, n1054);
  and g1834 (n1055, n_1041, n_1042);
  not g1843 (n_1043, n1063);
  and g1844 (n1064, n1055, n_1043);
  not g1845 (n_1044, n1044);
  and g1846 (n1065, n_1044, n1063);
  not g1847 (n_1045, n1064);
  not g1848 (n_1046, n1065);
  and g1849 (n1066, n_1045, n_1046);
  not g1858 (n_1047, n1074);
  and g1859 (n1075, n1066, n_1047);
  not g1860 (n_1048, n1055);
  and g1861 (n1076, n_1048, n1074);
  or g1862 (\P[4] , n1075, n1076);
  and g1863 (n1078, n1009, n1014);
  not g1889 (n_1049, n1103);
  and g1890 (n1104, n1087, n_1049);
  not g1891 (n_1050, n1078);
  or g1892 (\P[5] , n_1050, n1104);
  not g1893 (n_1051, n1087);
  or g1894 (\P[6] , n_1050, n_1051);
  and g1909 (n1005, n_583, n_570, n896, n744);
  and g1911 (n998, n_543, n_530, n886, n728);
  and g1913 (n991, n_503, n_490, n876, n712);
  and g1915 (n984, n_463, n_450, n866, n696);
  and g1917 (n977, n_423, n_410, n856, n680);
  and g1919 (n970, n_383, n_370, n846, n664);
  and g1921 (n963, n_343, n_330, n836, n648);
  and g1923 (n956, n_303, n_290, n826, n632);
  and g1925 (n949, n_263, n_250, n816, n616);
  and g1927 (n942, n_223, n_210, n806, n600);
  and g1929 (n935, n_183, n_170, n796, n584);
  and g1933 (n925, n_123, n568, n564, n560);
  and g1934 (n913, n_60, n532, n_73, n764);
  and g1936 (n917, n_103, n_90, n776, n552);
  and g1937 (n_1081, n_553, n_540, n_543);
  and g1938 (n_1082, n_530, n_533);
  and g1939 (n_1083, n_520, n_523);
  and g1940 (n_1084, n_510, n991);
  and g1941 (n1074, n_1081, n_1082, n_1083, n_1084);
  and g1942 (n_1085, n_473, n_460, n_463);
  and g1943 (n_1086, n_450, n_453);
  and g1944 (n_1087, n_440, n_443);
  and g1945 (n_1088, n_430, n977);
  and g1946 (n1063, n_1085, n_1086, n_1087, n_1088);
  and g1947 (n_1089, n_393, n_380, n_383);
  and g1948 (n_1090, n_370, n_373);
  and g1949 (n_1091, n_360, n_363);
  and g1950 (n_1092, n_350, n963);
  and g1951 (n1052, n_1089, n_1090, n_1091, n_1092);
  and g1952 (n_1093, n_313, n_300, n_303, n_290);
  and g1953 (n_1094, n_293, n_280, n_283, n_270);
  and g1954 (n_1095, n_273, n_260, n_263, n_250);
  and g1955 (n_1096, n_253, n_240, n_243);
  and g1956 (n1038, n_1093, n_1094, n_1095, n_1096);
  and g1957 (n_1097, n_130, n786);
  and g1959 (n1014, n_143, n917, n_1097, n568);
  and g1960 (n_1099, n_233, n_220, n_223);
  and g1961 (n_1100, n_210, n_213);
  and g1962 (n_1101, n_200, n_203);
  and g1963 (n_1102, n_190, n935);
  and g1964 (n1022, n_1099, n_1100, n_1101, n_1102);
  and g1965 (n_1103, n_270, n949, n_313);
  and g1966 (n_1104, n_300, n_303, n_290);
  and g1968 (n_1106, n_283, n1022);
  and g1969 (n1087, n_1103, n_1104, n624, n_1106);
  and g1971 (n_1108, n_463, n_450, n_453, n_440);
  and g1972 (n_1109, n_443, n_430, n_433, n_420);
  and g1973 (n_1110, n_423, n_410, n_413, n_400);
  and g1974 (n_1111, n_403, n_390, n1052, n696);
  and g1975 (n1103, n_1108, n_1109, n_1110, n_1111);
  nand g1976 (n_1113, n_621, n_610, n1005);
  nand g1977 (n_1114, n906, n1074);
  or g1978 (n_1115, n_1049, \A[0] );
  or g1980 (n_1116, \P[6] , \A[1] );
  or g1981 (F, n_1113, n_1114, n_1115, n_1116);
endmodule

