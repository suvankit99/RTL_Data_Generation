
module bar(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] ,
     \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14]
     , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
     \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
     \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
     \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
     \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
     \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
     \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
     \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
     \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
     \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
     \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
     \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
     \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105]
     , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] ,
     \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
     \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
     \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
     \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
     \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
     \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
     \result[10] , \result[11] , \result[12] , \result[13] ,
     \result[14] , \result[15] , \result[16] , \result[17] ,
     \result[18] , \result[19] , \result[20] , \result[21] ,
     \result[22] , \result[23] , \result[24] , \result[25] ,
     \result[26] , \result[27] , \result[28] , \result[29] ,
     \result[30] , \result[31] , \result[32] , \result[33] ,
     \result[34] , \result[35] , \result[36] , \result[37] ,
     \result[38] , \result[39] , \result[40] , \result[41] ,
     \result[42] , \result[43] , \result[44] , \result[45] ,
     \result[46] , \result[47] , \result[48] , \result[49] ,
     \result[50] , \result[51] , \result[52] , \result[53] ,
     \result[54] , \result[55] , \result[56] , \result[57] ,
     \result[58] , \result[59] , \result[60] , \result[61] ,
     \result[62] , \result[63] , \result[64] , \result[65] ,
     \result[66] , \result[67] , \result[68] , \result[69] ,
     \result[70] , \result[71] , \result[72] , \result[73] ,
     \result[74] , \result[75] , \result[76] , \result[77] ,
     \result[78] , \result[79] , \result[80] , \result[81] ,
     \result[82] , \result[83] , \result[84] , \result[85] ,
     \result[86] , \result[87] , \result[88] , \result[89] ,
     \result[90] , \result[91] , \result[92] , \result[93] ,
     \result[94] , \result[95] , \result[96] , \result[97] ,
     \result[98] , \result[99] , \result[100] , \result[101] ,
     \result[102] , \result[103] , \result[104] , \result[105] ,
     \result[106] , \result[107] , \result[108] , \result[109] ,
     \result[110] , \result[111] , \result[112] , \result[113] ,
     \result[114] , \result[115] , \result[116] , \result[117] ,
     \result[118] , \result[119] , \result[120] , \result[121] ,
     \result[122] , \result[123] , \result[124] , \result[125] ,
     \result[126] , \result[127] );
  input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
       \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
       \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
       \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
       \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
       \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] ,
       \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
       \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
       \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] ,
       \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] ,
       \shift[1] , \shift[2] , \shift[3] , \shift[4] , \shift[5] ,
       \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4]
       , \result[5] , \result[6] , \result[7] , \result[8] , \result[9]
       , \result[10] , \result[11] , \result[12] , \result[13] ,
       \result[14] , \result[15] , \result[16] , \result[17] ,
       \result[18] , \result[19] , \result[20] , \result[21] ,
       \result[22] , \result[23] , \result[24] , \result[25] ,
       \result[26] , \result[27] , \result[28] , \result[29] ,
       \result[30] , \result[31] , \result[32] , \result[33] ,
       \result[34] , \result[35] , \result[36] , \result[37] ,
       \result[38] , \result[39] , \result[40] , \result[41] ,
       \result[42] , \result[43] , \result[44] , \result[45] ,
       \result[46] , \result[47] , \result[48] , \result[49] ,
       \result[50] , \result[51] , \result[52] , \result[53] ,
       \result[54] , \result[55] , \result[56] , \result[57] ,
       \result[58] , \result[59] , \result[60] , \result[61] ,
       \result[62] , \result[63] , \result[64] , \result[65] ,
       \result[66] , \result[67] , \result[68] , \result[69] ,
       \result[70] , \result[71] , \result[72] , \result[73] ,
       \result[74] , \result[75] , \result[76] , \result[77] ,
       \result[78] , \result[79] , \result[80] , \result[81] ,
       \result[82] , \result[83] , \result[84] , \result[85] ,
       \result[86] , \result[87] , \result[88] , \result[89] ,
       \result[90] , \result[91] , \result[92] , \result[93] ,
       \result[94] , \result[95] , \result[96] , \result[97] ,
       \result[98] , \result[99] , \result[100] , \result[101] ,
       \result[102] , \result[103] , \result[104] , \result[105] ,
       \result[106] , \result[107] , \result[108] , \result[109] ,
       \result[110] , \result[111] , \result[112] , \result[113] ,
       \result[114] , \result[115] , \result[116] , \result[117] ,
       \result[118] , \result[119] , \result[120] , \result[121] ,
       \result[122] , \result[123] , \result[124] , \result[125] ,
       \result[126] , \result[127] ;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
       \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
       \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
       \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
       \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
       \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] ,
       \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
       \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
       \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] ,
       \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] ,
       \shift[1] , \shift[2] , \shift[3] , \shift[4] , \shift[5] ,
       \shift[6] ;
  wire \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
       \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
       \result[10] , \result[11] , \result[12] , \result[13] ,
       \result[14] , \result[15] , \result[16] , \result[17] ,
       \result[18] , \result[19] , \result[20] , \result[21] ,
       \result[22] , \result[23] , \result[24] , \result[25] ,
       \result[26] , \result[27] , \result[28] , \result[29] ,
       \result[30] , \result[31] , \result[32] , \result[33] ,
       \result[34] , \result[35] , \result[36] , \result[37] ,
       \result[38] , \result[39] , \result[40] , \result[41] ,
       \result[42] , \result[43] , \result[44] , \result[45] ,
       \result[46] , \result[47] , \result[48] , \result[49] ,
       \result[50] , \result[51] , \result[52] , \result[53] ,
       \result[54] , \result[55] , \result[56] , \result[57] ,
       \result[58] , \result[59] , \result[60] , \result[61] ,
       \result[62] , \result[63] , \result[64] , \result[65] ,
       \result[66] , \result[67] , \result[68] , \result[69] ,
       \result[70] , \result[71] , \result[72] , \result[73] ,
       \result[74] , \result[75] , \result[76] , \result[77] ,
       \result[78] , \result[79] , \result[80] , \result[81] ,
       \result[82] , \result[83] , \result[84] , \result[85] ,
       \result[86] , \result[87] , \result[88] , \result[89] ,
       \result[90] , \result[91] , \result[92] , \result[93] ,
       \result[94] , \result[95] , \result[96] , \result[97] ,
       \result[98] , \result[99] , \result[100] , \result[101] ,
       \result[102] , \result[103] , \result[104] , \result[105] ,
       \result[106] , \result[107] , \result[108] , \result[109] ,
       \result[110] , \result[111] , \result[112] , \result[113] ,
       \result[114] , \result[115] , \result[116] , \result[117] ,
       \result[118] , \result[119] , \result[120] , \result[121] ,
       \result[122] , \result[123] , \result[124] , \result[125] ,
       \result[126] , \result[127] ;
  wire n264, n265, n266, n267, n269, n270, n271, n272;
  wire n274, n275, n276, n277, n278, n279, n280, n282;
  wire n283, n284, n285, n287, n288, n289, n291, n292;
  wire n293, n294, n296, n297, n298, n299, n301, n302;
  wire n303, n304, n305, n306, n307, n309, n310, n311;
  wire n312, n314, n315, n316, n318, n319, n320, n321;
  wire n322, n323, n324, n326, n327, n328, n329, n331;
  wire n332, n333, n334, n335, n336, n338, n339, n340;
  wire n341, n343, n344, n346, n347, n348, n349, n351;
  wire n352, n353, n354, n356, n357, n358, n359, n360;
  wire n361, n363, n364, n365, n366, n368, n369, n371;
  wire n372, n373, n375, n376, n377, n378, n380, n381;
  wire n382, n383, n385, n386, n387, n388, n389, n390;
  wire n392, n393, n394, n395, n397, n398, n400, n401;
  wire n402, n403, n405, n406, n407, n408, n410, n411;
  wire n412, n413, n414, n415, n417, n418, n419, n420;
  wire n422, n423, n425, n426, n427, n428, n429, n430;
  wire n431, n433, n434, n435, n436, n438, n439, n440;
  wire n441, n442, n443, n445, n446, n447, n448, n450;
  wire n451, n453, n454, n455, n456, n458, n459, n460;
  wire n461, n463, n464, n465, n466, n467, n468, n470;
  wire n471, n472, n473, n475, n476, n478, n479, n480;
  wire n482, n483, n484, n485, n486, n487, n489, n490;
  wire n491, n492, n494, n495, n496, n497, n498, n499;
  wire n501, n502, n503, n504, n506, n507, n509, n510;
  wire n511, n512, n514, n515, n516, n517, n519, n520;
  wire n521, n522, n523, n524, n526, n527, n528, n529;
  wire n531, n532, n534, n535, n536, n537, n538, n539;
  wire n541, n542, n543, n544, n546, n547, n548, n549;
  wire n550, n551, n553, n554, n555, n556, n558, n559;
  wire n561, n562, n563, n564, n566, n567, n568, n569;
  wire n571, n572, n573, n574, n575, n576, n578, n579;
  wire n580, n581, n583, n584, n586, n587, n589, n590;
  wire n591, n592, n594, n595, n596, n597, n599, n600;
  wire n601, n602, n603, n604, n606, n607, n608, n609;
  wire n611, n612, n614, n615, n616, n617, n619, n620;
  wire n621, n622, n624, n625, n626, n627, n628, n629;
  wire n631, n632, n633, n634, n636, n637, n639, n640;
  wire n641, n642, n643, n644, n646, n647, n648, n649;
  wire n651, n652, n653, n654, n655, n656, n658, n659;
  wire n660, n661, n663, n664, n666, n667, n668, n669;
  wire n671, n672, n673, n674, n676, n677, n678, n679;
  wire n680, n681, n683, n684, n685, n686, n688, n689;
  wire n691, n692, n694, n695, n697, n698, n699, n700;
  wire n702, n703, n704, n705, n707, n708, n709, n710;
  wire n711, n712, n714, n715, n716, n717, n719, n720;
  wire n722, n723, n724, n725, n727, n728, n729, n730;
  wire n732, n733, n734, n735, n736, n737, n739, n740;
  wire n741, n742, n744, n745, n747, n748, n749, n750;
  wire n751, n752, n754, n755, n756, n757, n759, n760;
  wire n761, n762, n763, n764, n766, n767, n768, n769;
  wire n771, n772, n774, n775, n776, n777, n779, n780;
  wire n781, n782, n784, n785, n786, n787, n788, n789;
  wire n791, n792, n793, n794, n796, n797, n799, n800;
  wire n802, n803, n804, n805, n807, n808, n809, n810;
  wire n812, n813, n814, n815, n816, n817, n819, n820;
  wire n821, n822, n824, n825, n827, n828, n829, n830;
  wire n832, n833, n834, n835, n837, n838, n839, n840;
  wire n841, n842, n844, n845, n846, n847, n849, n850;
  wire n852, n853, n854, n855, n856, n857, n859, n860;
  wire n861, n862, n864, n865, n866, n867, n868, n869;
  wire n871, n872, n873, n874, n876, n877, n879, n880;
  wire n881, n882, n884, n885, n886, n887, n889, n890;
  wire n891, n892, n893, n894, n896, n897, n898, n899;
  wire n901, n902, n904, n905, n907, n908, n909, n910;
  wire n911, n912, n914, n915, n916, n917, n919, n920;
  wire n921, n922, n923, n924, n926, n927, n928, n929;
  wire n931, n932, n934, n935, n936, n937, n939, n940;
  wire n941, n942, n944, n945, n946, n947, n948, n949;
  wire n951, n952, n953, n954, n956, n957, n959, n960;
  wire n961, n962, n963, n964, n966, n967, n968, n969;
  wire n971, n972, n973, n974, n975, n976, n978, n979;
  wire n980, n981, n983, n984, n986, n987, n988, n989;
  wire n991, n992, n993, n994, n996, n997, n998, n999;
  wire n1000, n1001, n1003, n1004, n1005, n1006, n1008, n1009;
  wire n1011, n1012, n1014, n1015, n1016, n1017, n1019, n1020;
  wire n1021, n1022, n1024, n1025, n1026, n1027, n1028, n1029;
  wire n1031, n1032, n1033, n1034, n1036, n1037, n1039, n1040;
  wire n1041, n1042, n1044, n1045, n1046, n1047, n1049, n1050;
  wire n1051, n1052, n1053, n1054, n1056, n1057, n1058, n1059;
  wire n1061, n1062, n1064, n1065, n1066, n1067, n1068, n1069;
  wire n1071, n1072, n1073, n1074, n1076, n1077, n1078, n1079;
  wire n1080, n1081, n1083, n1084, n1085, n1086, n1088, n1089;
  wire n1091, n1092, n1093, n1094, n1096, n1097, n1098, n1099;
  wire n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109;
  wire n1110, n1111, n1113, n1114, n1116, n1117, n1119, n1120;
  wire n1122, n1123, n1125, n1126, n1128, n1129, n1130, n1131;
  wire n1133, n1134, n1136, n1137, n1139, n1140, n1142, n1143;
  wire n1145, n1146, n1147, n1148, n1150, n1151, n1153, n1154;
  wire n1156, n1157, n1158, n1159, n1161, n1162, n1164, n1165;
  wire n1166, n1167, n1169, n1170, n1172, n1173, n1175, n1176;
  wire n1178, n1179, n1181, n1182, n1183, n1184, n1186, n1187;
  wire n1189, n1190, n1192, n1193, n1195, n1196, n1198, n1199;
  wire n1201, n1202, n1203, n1204, n1206, n1207, n1209, n1210;
  wire n1212, n1213, n1215, n1216, n1218, n1219, n1220, n1221;
  wire n1223, n1224, n1226, n1227, n1229, n1230, n1231, n1232;
  wire n1234, n1235, n1237, n1238, n1239, n1240, n1242, n1243;
  wire n1245, n1246, n1248, n1249, n1251, n1252, n1254, n1255;
  wire n1256, n1257, n1259, n1260, n1262, n1263, n1265, n1266;
  wire n1268, n1269, n1270, n1271, n1273, n1274, n1276, n1277;
  wire n1278, n1279, n1281, n1282, n1284, n1285, n1287, n1288;
  wire n1290, n1291, n1293, n1294, n1295, n1296, n1298, n1299;
  wire n1301, n1302, n1304, n1305, n1306, n1307, n1309, n1310;
  wire n1312, n1313, n1314, n1315, n1317, n1318, n1320, n1321;
  wire n1323, n1324, n1326, n1327, n1329, n1330, n1331, n1332;
  wire n1334, n1335, n1337, n1338, n1340, n1341, n1343, n1344;
  wire n1346, n1347, n1349, n1350, n1351, n1352, n1354, n1355;
  wire n1357, n1358, n1360, n1361, n1363, n1364, n1366, n1367;
  wire n1368, n1369, n1371, n1372, n1374, n1375, n1377, n1378;
  wire n1379, n1380, n1382, n1383, n1385, n1386, n1387, n1388;
  wire n1390, n1391, n1393, n1394, n1396, n1397, n1399, n1400;
  wire n1402, n1403, n1404, n1405, n1407, n1408, n1410, n1411;
  wire n1413, n1414, n1416, n1417, n1419, n1420, n1422, n1423;
  wire n1425, n1426, n1427, n1428, n1430, n1431, n1433, n1434;
  wire n1436, n1437, n1439, n1440, n1442, n1443, n1444, n1445;
  wire n1447, n1448, n1450, n1451, n1453, n1454, n1455, n1456;
  wire n1458, n1459, n1461, n1462, n1463, n1464, n1466, n1467;
  wire n1469, n1470, n1472, n1473, n1475, n1476, n1478, n1479;
  wire n1480, n1481, n1483, n1484, n1486, n1487, n1489, n1490;
  wire n1492, n1493, n1495, n1496, n1498, n1499, n1500, n1501;
  wire n1503, n1504, n1506, n1507, n1509, n1510, n1512, n1513;
  wire n1515, n1516, n1517, n1518, n1520, n1521, n1523, n1524;
  wire n1526, n1527, n1528, n1529, n1531, n1532, n1534, n1535;
  wire n1536, n1537, n1539, n1540, n1542, n1543, n1545, n1546;
  wire n1548, n1549, n1551, n1552, n1553, n1554, n1556, n1557;
  wire n1559, n1560, n1562, n1563, n1565, n1566, n1567, n1568;
  wire n1570, n1571, n1573, n1574, n1575, n1576, n1578, n1579;
  wire n1581, n1582, n1584, n1585, n1587, n1588, n1590, n1591;
  wire n1592, n1593, n1595, n1596, n1598, n1599, n1601, n1602;
  wire n1603, n1604, n1606, n1607, n1609, n1610, n1611, n1612;
  wire n1614, n1615, n1617, n1618, n1620, n1621, n1623, n1624;
  wire n1626, n1627, n1628, n1629, n1631, n1632, n1634, n1635;
  wire n1637, n1638, n1640, n1641, n1643, n1644, n1646, n1647;
  wire n1648, n1649, n1651, n1652, n1654, n1655, n1657, n1658;
  wire n1660, n1661, n1663, n1664, n1665, n1666, n1668, n1669;
  wire n1671, n1672, n1674, n1675, n1676, n1677, n1679, n1680;
  wire n1682, n1683, n1684, n1685, n1687, n1688, n1690, n1691;
  wire n1693, n1694, n1696, n1697, n1699, n1700, n1701, n1702;
  wire n1704, n1705, n1707, n1708, n1710, n1711, n1713, n1714;
  wire n1716, n1717, n1719, n1720, n1722, n1723, n1724, n1725;
  wire n1727, n1728, n1730, n1731, n1733, n1734, n1736, n1737;
  wire n1739, n1740, n1741, n1742, n1744, n1745, n1747, n1748;
  wire n1750, n1751, n1752, n1753, n1755, n1756, n1758, n1759;
  wire n1760, n1761, n1763, n1764, n1766, n1767, n1769, n1770;
  wire n1772, n1773, n1775, n1776, n1777, n1778, n1780, n1781;
  wire n1783, n1784, n1786, n1787, n1789, n1790, n1792, n1793;
  wire n1795, n1796, n1797, n1798, n1800, n1801, n1803, n1804;
  wire n1806, n1807, n1809, n1810, n1812, n1813, n1814, n1815;
  wire n1817, n1818, n1820, n1821, n1823, n1824, n1825, n1826;
  wire n1828, n1829, n1831, n1832, n1833, n1834, n1836, n1837;
  wire n1839, n1840, n1842, n1843, n1845, n1846, n1848, n1849;
  wire n1850, n1851, n1853, n1854, n1856, n1857, n1859, n1860;
  wire n1862, n1863, n1865, n1866, n1868, n1869, n1870, n1871;
  wire n1873, n1874, n1876, n1877, n1879, n1880, n1882, n1883;
  wire n1885, n1886, n1887, n1888, n1890, n1891, n1893, n1894;
  wire n1896, n1897, n1898, n1899, n1901, n1902, n1904, n1905;
  wire n1906, n1907, n1909, n1910, n1912, n1913, n1915, n1916;
  wire n1918, n1919, n1921, n1922, n1923, n1924, n1926, n1927;
  wire n1929, n1930, n1932, n1933, n1935, n1936, n1938, n1939;
  wire n1941, n1942, n1943, n1944, n1946, n1947, n1949, n1950;
  wire n1952, n1953, n1955, n1956, n1958, n1959, n1960, n1961;
  wire n1963, n1964, n1966, n1967, n1969, n1970, n1971, n1972;
  wire n1974, n1975, n1977, n1978, n1979, n1980, n1982, n1983;
  wire n1985, n1986, n1988, n1989, n1991, n1992, n1994, n1995;
  wire n1996, n1997, n1999, n2000, n2002, n2003, n2005, n2006;
  wire n2008, n2009, n2011, n2012, n2014, n2015, n2016, n2017;
  wire n2019, n2020, n2022, n2023, n2025, n2026, n2028, n2029;
  wire n2031, n2032, n2033, n2034, n2036, n2037, n2039, n2040;
  wire n2042, n2043, n2044, n2045, n2047, n2048, n2050, n2051;
  wire n2052, n2053, n2055, n2056, n2058, n2059, n2061, n2062;
  wire n2064, n2065, n2067, n2068, n2069, n2070, n2072, n2073;
  wire n2075, n2076, n2078, n2079, n2081, n2082, n2084, n2085;
  wire n2087, n2088, n2089, n2090, n2092, n2093, n2095, n2096;
  wire n2098, n2099, n2101, n2102, n2104, n2105, n2106, n2107;
  wire n2109, n2110, n2112, n2113, n2115, n2116, n2117, n2118;
  wire n2120, n2121, n2123, n2124, n2125, n2126, n2128, n2129;
  wire n2131, n2132, n2134, n2135, n2137, n2138, n2140, n2141;
  wire n2142, n2143, n2145, n2146, n2148, n2149, n2151, n2152;
  wire n2154, n2155, n2157, n2158, n2160, n2161, n2162, n2163;
  wire n2165, n2166, n2168, n2169, n2171, n2172, n2174, n2175;
  wire n2177, n2178, n2179, n2180, n2182, n2183, n2185, n2186;
  wire n2188, n2189, n2190, n2191, n2193, n2194, n2196, n2197;
  wire n2198, n2199, n2201, n2202, n2204, n2205, n2207, n2208;
  wire n2210, n2211, n2213, n2214, n2215, n2216, n2218, n2219;
  wire n2221, n2222, n2224, n2225, n2227, n2228, n2230, n2231;
  wire n2233, n2234, n2235, n2236, n2238, n2239, n2241, n2242;
  wire n2244, n2245, n2247, n2248, n2250, n2251, n2252, n2253;
  wire n2255, n2256, n2258, n2259, n2261, n2262, n2263, n2264;
  wire n2266, n2267, n2269, n2270, n2271, n2272, n2274, n2275;
  wire n2277, n2278, n2280, n2281, n2283, n2284, n2286, n2287;
  wire n2288, n2289, n2291, n2292, n2294, n2295, n2297, n2298;
  wire n2300, n2301, n2303, n2304, n2306, n2307, n2308, n2309;
  wire n2311, n2312, n2314, n2315, n2317, n2318, n2320, n2321;
  wire n2323, n2324, n2325, n2326, n2328, n2329, n2331, n2332;
  wire n2334, n2335, n2336, n2337, n2339, n2340, n2342, n2343;
  wire n2344, n2345, n2347, n2348, n2350, n2351, n2353, n2354;
  wire n2356, n2357, n2359, n2360, n2361, n2362, n2364, n2365;
  wire n2367, n2368, n2370, n2371, n2373, n2374, n2376, n2377;
  wire n2379, n2380, n2381, n2382, n2384, n2385, n2387, n2388;
  wire n2390, n2391, n2393, n2394, n2396, n2397, n2398, n2399;
  wire n2401, n2402, n2404, n2405, n2407, n2408, n2409, n2410;
  wire n2412, n2413, n2415, n2416, n2417, n2418, n2420, n2421;
  wire n2423, n2424, n2426, n2427, n2429, n2430, n2432, n2433;
  wire n2434, n2435, n2437, n2438, n2440, n2441, n2443, n2444;
  wire n2446, n2447, n2449, n2450, n2452, n2453, n2454, n2455;
  wire n2457, n2458, n2460, n2461, n2463, n2464, n2466, n2467;
  wire n2469, n2470, n2471, n2472, n2474, n2475, n2477, n2478;
  wire n2480, n2481, n2482, n2483, n2485, n2486, n2488, n2489;
  wire n2490, n2491, n2493, n2494, n2496, n2497, n2499, n2500;
  wire n2502, n2503, n2505, n2506, n2507, n2508, n2510, n2511;
  wire n2513, n2514, n2516, n2517, n2519, n2520, n2522, n2523;
  wire n2525, n2526, n2527, n2528, n2530, n2531, n2533, n2534;
  wire n2536, n2537, n2539, n2540, n2542, n2543, n2544, n2545;
  wire n2547, n2548, n2550, n2551, n2553, n2554, n2555, n2556;
  wire n2558, n2559, n2561, n2562, n2563, n2564, n2566, n2567;
  wire n2569, n2570, n2572, n2573, n2575, n2576, n2578, n2579;
  wire n2580, n2581, n2583, n2584, n2586, n2587, n2589, n2590;
  wire n2592, n2593, n2595, n2596, n2598, n2599, n2600, n2601;
  wire n2603, n2604, n2606, n2607, n2609, n2610, n2612, n2613;
  wire n2615, n2616, n2617, n2618, n2620, n2621, n2623, n2624;
  wire n2626, n2627, n2629, n2630, n2632, n2633, n2634, n2635;
  wire n2637, n2638, n2640, n2641, n2643, n2644, n2646, n2647;
  wire n2649, n2650, n2651, n2652, n2654, n2655, n2657, n2658;
  wire n2660, n2661, n2663, n2664, n2666, n2667, n2668, n2669;
  wire n2671, n2672, n2674, n2675, n2677, n2678, n2680, n2681;
  wire n2683, n2684, n2685, n2686, n2688, n2689, n2691, n2692;
  wire n2694, n2695, n2697, n2698, n2700, n2701, n2702, n2703;
  wire n2705, n2706, n2708, n2709, n2711, n2712, n2714, n2715;
  wire n2717, n2718, n2719, n2720, n2722, n2723, n2725, n2726;
  wire n2728, n2729, n2731, n2732, n2734, n2735, n2736, n2737;
  wire n2739, n2740, n2742, n2743, n2745, n2746, n2748, n2749;
  wire n2751, n2752, n2753, n2754, n2756, n2757, n2759, n2760;
  wire n2762, n2763, n2765, n2766, n2768, n2769, n2770, n2771;
  wire n2773, n2774, n2776, n2777, n2779, n2780, n2782, n2783;
  wire n2785, n2786, n2787, n2788, n2790, n2791, n2793, n2794;
  wire n2796, n2797, n2799, n2800, n2802, n2803, n2804, n2805;
  wire n2807, n2808, n2810, n2811, n2813, n2814, n2816, n2817;
  wire n2819, n2820, n2821, n2822, n2824, n2825, n2827, n2828;
  wire n2830, n2831, n2833, n2834, n2836, n2837, n2838, n2839;
  wire n2841, n2842, n2844, n2845, n2847, n2848, n2850, n2851;
  wire n2853, n2854, n2855, n2856, n2858, n2859, n2861, n2862;
  wire n2864, n2865, n2867, n2868, n2870, n2871, n2872, n2873;
  wire n2875, n2876, n2878, n2879, n2881, n2882, n2884, n2885;
  wire n2887, n2888, n2889, n2890, n2892, n2893, n2895, n2896;
  wire n2898, n2899, n2901, n2902, n2904, n2905, n2906, n2907;
  wire n2909, n2910, n2912, n2913, n2915, n2916, n2918, n2919;
  wire n2921, n2922, n2923, n2924, n2926, n2927, n2929, n2930;
  wire n2932, n2933, n2935, n2936, n2938, n2939, n2940, n2941;
  wire n2943, n2944, n2946, n2947, n2949, n2950, n2952, n2953;
  wire n2955, n2956, n2957, n2958, n2960, n2961, n2963, n2964;
  wire n2966, n2967, n2969, n2970, n2972, n2973, n2974, n2975;
  wire n2977, n2978, n2980, n2981, n2983, n2984, n2986, n2987;
  wire n2989, n2990, n2991, n2992, n2994, n2995, n2997, n2998;
  wire n3000, n3001, n3003, n3004, n3006, n3007, n3008, n3009;
  wire n3011, n3012, n3014, n3015, n3017, n3018, n3020, n3021;
  wire n3023, n3024, n3025, n3026, n3028, n3029, n3031, n3032;
  wire n3034, n3035, n3037, n3038, n3040, n3041, n3042, n3043;
  wire n3045, n3046, n3048, n3049, n3051, n3052, n3054, n3055;
  wire n3057, n3058, n3059, n3060, n3062, n3063, n3065, n3066;
  wire n3068, n3069, n3071, n3072, n3074, n3075, n3076, n3077;
  wire n3079, n3080, n3082, n3083, n3085, n3086, n3088, n3089;
  wire n3091, n3092, n3093, n3094, n3096, n3097, n3099, n3100;
  wire n3102, n3103, n3105, n3106, n3108, n3109, n3110, n3111;
  wire n3113, n3114, n3116, n3117, n3119, n3120, n3122, n3123;
  wire n3125, n3126, n3127, n3128, n3130, n3131, n3133, n3134;
  wire n3136, n3137, n3139, n3140, n3142, n3143, n3144, n3145;
  wire n3147, n3148, n3150, n3151, n3153, n3154, n3156, n3157;
  wire n3159, n3160, n3161, n3162, n3164, n3165, n3167, n3168;
  wire n3170, n3171, n3173, n3174, n3176, n3177, n3178, n3179;
  wire n3181, n3182, n3184, n3185, n3187, n3188, n3190, n3191;
  wire n3193, n3194, n3195, n3196, n3198, n3199, n3201, n3202;
  wire n3204, n3205, n3207, n3208, n3210, n3211, n3212, n3213;
  wire n3215, n3216, n3218, n3219, n3221, n3222, n3224, n3225;
  wire n3227, n3228, n3229, n3230, n3232, n3233, n3235, n3236;
  wire n3238, n3239, n3241, n3242, n3244, n3245, n3246, n3247;
  wire n3249, n3250, n3252, n3253, n3255, n3256, n3258, n3259;
  wire n3261, n3262, n3263, n3264, n3266, n3267, n3269, n3270;
  wire n3272, n3273, n3275, n3276, n3278, n3279, n3280, n3281;
  wire n3283, n3284, n3286, n3287, n3289, n3290, n3292, n3293;
  wire n3295, n3296, n3297, n3298, n3300, n3301, n3303, n3304;
  wire n3306, n3307, n3309, n3310, n3312, n3313, n3314, n3315;
  wire n3317, n3318, n3320, n3321, n3323, n3324, n3326, n3327;
  wire n3329, n3330, n3331, n3332, n3334, n3335, n3337, n3338;
  wire n3340, n3341, n3343, n3344, n3346, n3347, n3348, n3349;
  wire n3351, n3352, n3354, n3355, n3357, n3358, n3360, n3361;
  wire n3363, n3364, n3365, n3366, n3368, n3369, n3371, n3372;
  wire n3374, n3375, n3377, n3378, n3380, n3381, n3382, n3383;
  wire n3385, n3386, n3388, n3389, n3391, n3392, n3394, n3395;
  wire n3397, n3398, n3399, n3400, n3402, n3403, n3405, n3406;
  wire n3408, n3409, n3411, n3412, n3414, n3415, n3417, n3418;
  wire n3420, n3421, n3423, n3424, n3426, n3427, n3429, n3430;
  wire n3432, n3433, n3435, n3436, n3438, n3439, n3441, n3442;
  wire n3444, n3445, n3447, n3448, n3450, n3451, n3453, n3454;
  wire n3456, n3457, n3459, n3460, n3462, n3463, n3465, n3466;
  wire n3468, n3469, n3471, n3472, n3474, n3475, n3477, n3478;
  wire n3480, n3481, n3483, n3484, n3486, n3487, n3489, n3490;
  wire n3492, n3493, n3495, n3496, n3498, n3499, n3501, n3502;
  wire n3504, n3505, n3507, n3508, n3510, n3511, n3513, n3514;
  wire n3516, n3517, n3519, n3520, n3522, n3523, n3525, n3526;
  wire n3528, n3529, n3531, n3532, n3534, n3535, n3537, n3538;
  wire n3540, n3541, n3543, n3544, n3546, n3547, n3549, n3550;
  wire n3552, n3553, n3555, n3556, n3558, n3559, n3561, n3562;
  wire n3564, n3565, n3567, n3568, n3570, n3571, n3573, n3574;
  wire n3576, n3577, n3579, n3580, n3582, n3583, n3585, n3586;
  wire n3588, n3589, n3591, n3592, n3594, n3595, n3597, n3598;
  wire n_5, n_9, n_15, n_16, n_17, n_26, n_37, n_46;
  wire n_51, n_60, n_69, n_80, n_89, n_92, n_93, n_104;
  wire n_113, n_124, n_133, n_136, n_137, n_146, n_155, n_166;
  wire n_175, n_178, n_182, n_183, n_192, n_201, n_212, n_221;
  wire n_224, n_233, n_242, n_253, n_262, n_265, n_276, n_285;
  wire n_296, n_305, n_308, n_317, n_326, n_337, n_346, n_349;
  wire n_352, n_357, n_362, n_369, n_374, n_377, n_382, n_387;
  wire n_394, n_399, n_402, n_409, n_414, n_421, n_426, n_429;
  wire n_434, n_439, n_446, n_451, n_454, n_457, n_462, n_467;
  wire n_474, n_479, n_482, n_487, n_492, n_499, n_504, n_507;
  wire n_514, n_519, n_526, n_531, n_534, n_539, n_544, n_551;
  wire n_556, n_559, n_562, n_567, n_572, n_579, n_584, n_587;
  wire n_592, n_597, n_604, n_609, n_612, n_619, n_624, n_631;
  wire n_636, n_639, n_644, n_649, n_656, n_661, n_664, n_667;
  wire n_672, n_677, n_684, n_689, n_692, n_697, n_702, n_709;
  wire n_714, n_717, n_724, n_729, n_736, n_741, n_744, n_749;
  wire n_754, n_761, n_766, n_769, n_772, n_777, n_782, n_789;
  wire n_794, n_797, n_802, n_807, n_814, n_819, n_822, n_829;
  wire n_834, n_841, n_846, n_849, n_854, n_859, n_866, n_871;
  wire n_874, n_877, n_882, n_887, n_894, n_899, n_902, n_907;
  wire n_912, n_919, n_924, n_927, n_934, n_939, n_946, n_951;
  wire n_954, n_959, n_964, n_971, n_976, n_979, n_982, n_987;
  wire n_992, n_999, n_1004, n_1007, n_1012, n_1017, n_1024, n_1029;
  wire n_1032, n_1037, n_1042, n_1049, n_1054, n_1057, n_1062, n_1067;
  wire n_1074, n_1079, n_1082, n_1087, n_1092, n_1099, n_1104, n_1107;
  wire n_1112, n_1117, n_1124, n_1129, n_1132, n_1137, n_1142, n_1149;
  wire n_1154, n_1157, n_1162, n_1167, n_1174, n_1179, n_1182, n_1187;
  wire n_1192, n_1199, n_1204, n_1207, n_1212, n_1217, n_1224, n_1229;
  wire n_1232, n_1237, n_1242, n_1249, n_1254, n_1257, n_1262, n_1267;
  wire n_1274, n_1279, n_1282, n_1287, n_1292, n_1299, n_1304, n_1307;
  wire n_1312, n_1317, n_1324, n_1329, n_1332, n_1337, n_1342, n_1349;
  wire n_1354, n_1357, n_1362, n_1367, n_1374, n_1379, n_1382, n_1387;
  wire n_1392, n_1399, n_1404, n_1407, n_1412, n_1417, n_1424, n_1429;
  wire n_1432, n_1437, n_1442, n_1449, n_1454, n_1457, n_1462, n_1467;
  wire n_1474, n_1479, n_1482, n_1487, n_1492, n_1499, n_1504, n_1507;
  wire n_1512, n_1517, n_1524, n_1529, n_1532, n_1537, n_1542, n_1549;
  wire n_1554, n_1557, n_1562, n_1567, n_1574, n_1579, n_1582, n_1587;
  wire n_1592, n_1597, n_1602, n_1607, n_1612, n_1617, n_1622, n_1627;
  wire n_1632, n_1637, n_1642, n_1647, n_1652, n_1657, n_1662, n_1667;
  wire n_1672, n_1677, n_1682, n_1687, n_1692, n_1697, n_1702, n_1707;
  wire n_1712, n_1717, n_1722, n_1727, n_1732, n_1737, n_1742, n_1747;
  wire n_1752, n_1757, n_1762, n_1767, n_1772, n_1777, n_1782, n_1787;
  wire n_1792, n_1797, n_1802, n_1807, n_1812, n_1817, n_1822, n_1827;
  wire n_1832, n_1837, n_1842, n_1847, n_1852, n_1857, n_1862, n_1867;
  wire n_1872, n_1877, n_1882, n_1887, n_1892, n_1897, n_1902, n_1907;
  wire n_1912, n_1917, n_1922, n_1927, n_1932, n_1937, n_1942, n_1947;
  wire n_1952, n_1957, n_1962, n_1967, n_1972, n_1977, n_1982, n_1987;
  wire n_1992, n_1997, n_2002, n_2007, n_2012, n_2017, n_2022, n_2027;
  wire n_2032, n_2037, n_2042, n_2047, n_2052, n_2057, n_2062;
  and g1 (n264, \a[77] , \shift[0] );
  and g2 (n265, \shift[1] , n264);
  not g3 (n_5, \shift[0] );
  and g4 (n266, \a[78] , n_5);
  and g5 (n267, \shift[1] , n266);
  and g9 (n269, \a[80] , n_5);
  not g10 (n_9, \shift[1] );
  and g11 (n270, n_9, n269);
  and g12 (n271, \a[79] , \shift[0] );
  and g13 (n272, n_9, n271);
  not g18 (n_15, \shift[2] );
  not g19 (n_16, \shift[3] );
  and g20 (n275, n_15, n_16);
  not g21 (n_17, n274);
  and g22 (n276, n_17, n275);
  and g23 (n277, \a[73] , \shift[0] );
  and g24 (n278, \shift[1] , n277);
  and g25 (n279, \a[74] , n_5);
  and g26 (n280, \shift[1] , n279);
  and g30 (n282, \a[76] , n_5);
  and g31 (n283, n_9, n282);
  and g32 (n284, \a[75] , \shift[0] );
  and g33 (n285, n_9, n284);
  and g38 (n288, \shift[2] , n_16);
  not g39 (n_26, n287);
  and g40 (n289, n_26, n288);
  and g44 (n291, \a[65] , \shift[0] );
  and g45 (n292, \shift[1] , n291);
  and g46 (n293, \a[66] , n_5);
  and g47 (n294, \shift[1] , n293);
  and g51 (n296, \a[68] , n_5);
  and g52 (n297, n_9, n296);
  and g53 (n298, \a[67] , \shift[0] );
  and g54 (n299, n_9, n298);
  and g59 (n302, \shift[2] , \shift[3] );
  not g60 (n_37, n301);
  and g61 (n303, n_37, n302);
  and g62 (n304, \a[69] , \shift[0] );
  and g63 (n305, \shift[1] , n304);
  and g64 (n306, \a[70] , n_5);
  and g65 (n307, \shift[1] , n306);
  and g69 (n309, \a[72] , n_5);
  and g70 (n310, n_9, n309);
  and g71 (n311, \a[71] , \shift[0] );
  and g72 (n312, n_9, n311);
  and g77 (n315, n_15, \shift[3] );
  not g78 (n_46, n314);
  and g79 (n316, n_46, n315);
  and g84 (n319, \shift[4] , \shift[5] );
  not g85 (n_51, n318);
  and g86 (n320, n_51, n319);
  and g87 (n321, \a[93] , \shift[0] );
  and g88 (n322, \shift[1] , n321);
  and g89 (n323, \a[94] , n_5);
  and g90 (n324, \shift[1] , n323);
  and g94 (n326, \a[96] , n_5);
  and g95 (n327, n_9, n326);
  and g96 (n328, \a[95] , \shift[0] );
  and g97 (n329, n_9, n328);
  not g102 (n_60, n331);
  and g103 (n332, n275, n_60);
  and g104 (n333, \a[89] , \shift[0] );
  and g105 (n334, \shift[1] , n333);
  and g106 (n335, \a[90] , n_5);
  and g107 (n336, \shift[1] , n335);
  and g111 (n338, \a[92] , n_5);
  and g112 (n339, n_9, n338);
  and g113 (n340, \a[91] , \shift[0] );
  and g114 (n341, n_9, n340);
  not g119 (n_69, n343);
  and g120 (n344, n288, n_69);
  and g124 (n346, \a[81] , \shift[0] );
  and g125 (n347, \shift[1] , n346);
  and g126 (n348, \a[82] , n_5);
  and g127 (n349, \shift[1] , n348);
  and g131 (n351, \a[84] , n_5);
  and g132 (n352, n_9, n351);
  and g133 (n353, \a[83] , \shift[0] );
  and g134 (n354, n_9, n353);
  not g139 (n_80, n356);
  and g140 (n357, n302, n_80);
  and g141 (n358, \a[85] , \shift[0] );
  and g142 (n359, \shift[1] , n358);
  and g143 (n360, \a[86] , n_5);
  and g144 (n361, \shift[1] , n360);
  and g148 (n363, \a[88] , n_5);
  and g149 (n364, n_9, n363);
  and g150 (n365, \a[87] , \shift[0] );
  and g151 (n366, n_9, n365);
  not g156 (n_89, n368);
  and g157 (n369, n315, n_89);
  not g162 (n_92, \shift[4] );
  and g163 (n372, n_92, \shift[5] );
  not g164 (n_93, n371);
  and g165 (n373, n_93, n372);
  and g169 (n375, \a[125] , \shift[0] );
  and g170 (n376, \shift[1] , n375);
  and g171 (n377, \a[126] , n_5);
  and g172 (n378, \shift[1] , n377);
  and g176 (n380, \a[0] , n_5);
  and g177 (n381, n_9, n380);
  and g178 (n382, \a[127] , \shift[0] );
  and g179 (n383, n_9, n382);
  not g184 (n_104, n385);
  and g185 (n386, n275, n_104);
  and g186 (n387, \a[121] , \shift[0] );
  and g187 (n388, \shift[1] , n387);
  and g188 (n389, \a[122] , n_5);
  and g189 (n390, \shift[1] , n389);
  and g193 (n392, \a[124] , n_5);
  and g194 (n393, n_9, n392);
  and g195 (n394, \a[123] , \shift[0] );
  and g196 (n395, n_9, n394);
  not g201 (n_113, n397);
  and g202 (n398, n288, n_113);
  and g206 (n400, \a[113] , \shift[0] );
  and g207 (n401, \shift[1] , n400);
  and g208 (n402, \a[114] , n_5);
  and g209 (n403, \shift[1] , n402);
  and g213 (n405, \a[116] , n_5);
  and g214 (n406, n_9, n405);
  and g215 (n407, \a[115] , \shift[0] );
  and g216 (n408, n_9, n407);
  not g221 (n_124, n410);
  and g222 (n411, n302, n_124);
  and g223 (n412, \a[117] , \shift[0] );
  and g224 (n413, \shift[1] , n412);
  and g225 (n414, \a[118] , n_5);
  and g226 (n415, \shift[1] , n414);
  and g230 (n417, \a[120] , n_5);
  and g231 (n418, n_9, n417);
  and g232 (n419, \a[119] , \shift[0] );
  and g233 (n420, n_9, n419);
  not g238 (n_133, n422);
  and g239 (n423, n315, n_133);
  not g244 (n_136, \shift[5] );
  and g245 (n426, n_92, n_136);
  not g246 (n_137, n425);
  and g247 (n427, n_137, n426);
  and g248 (n428, \a[109] , \shift[0] );
  and g249 (n429, \shift[1] , n428);
  and g250 (n430, \a[110] , n_5);
  and g251 (n431, \shift[1] , n430);
  and g255 (n433, \a[112] , n_5);
  and g256 (n434, n_9, n433);
  and g257 (n435, \a[111] , \shift[0] );
  and g258 (n436, n_9, n435);
  not g263 (n_146, n438);
  and g264 (n439, n275, n_146);
  and g265 (n440, \a[105] , \shift[0] );
  and g266 (n441, \shift[1] , n440);
  and g267 (n442, \a[106] , n_5);
  and g268 (n443, \shift[1] , n442);
  and g272 (n445, \a[108] , n_5);
  and g273 (n446, n_9, n445);
  and g274 (n447, \a[107] , \shift[0] );
  and g275 (n448, n_9, n447);
  not g280 (n_155, n450);
  and g281 (n451, n288, n_155);
  and g285 (n453, \a[97] , \shift[0] );
  and g286 (n454, \shift[1] , n453);
  and g287 (n455, \a[98] , n_5);
  and g288 (n456, \shift[1] , n455);
  and g292 (n458, \a[100] , n_5);
  and g293 (n459, n_9, n458);
  and g294 (n460, \a[99] , \shift[0] );
  and g295 (n461, n_9, n460);
  not g300 (n_166, n463);
  and g301 (n464, n302, n_166);
  and g302 (n465, \a[101] , \shift[0] );
  and g303 (n466, \shift[1] , n465);
  and g304 (n467, \a[102] , n_5);
  and g305 (n468, \shift[1] , n467);
  and g309 (n470, \a[104] , n_5);
  and g310 (n471, n_9, n470);
  and g311 (n472, \a[103] , \shift[0] );
  and g312 (n473, n_9, n472);
  not g317 (n_175, n475);
  and g318 (n476, n315, n_175);
  and g323 (n479, \shift[4] , n_136);
  not g324 (n_178, n478);
  and g325 (n480, n_178, n479);
  not g330 (n_182, \shift[6] );
  not g331 (n_183, n482);
  and g332 (n483, n_182, n_183);
  and g333 (n484, \a[13] , \shift[0] );
  and g334 (n485, \shift[1] , n484);
  and g335 (n486, \a[14] , n_5);
  and g336 (n487, \shift[1] , n486);
  and g340 (n489, \a[16] , n_5);
  and g341 (n490, n_9, n489);
  and g342 (n491, \a[15] , \shift[0] );
  and g343 (n492, n_9, n491);
  not g348 (n_192, n494);
  and g349 (n495, n275, n_192);
  and g350 (n496, \a[9] , \shift[0] );
  and g351 (n497, \shift[1] , n496);
  and g352 (n498, \a[10] , n_5);
  and g353 (n499, \shift[1] , n498);
  and g357 (n501, \a[12] , n_5);
  and g358 (n502, n_9, n501);
  and g359 (n503, \a[11] , \shift[0] );
  and g360 (n504, n_9, n503);
  not g365 (n_201, n506);
  and g366 (n507, n288, n_201);
  and g370 (n509, \a[1] , \shift[0] );
  and g371 (n510, \shift[1] , n509);
  and g372 (n511, \a[2] , n_5);
  and g373 (n512, \shift[1] , n511);
  and g377 (n514, \a[4] , n_5);
  and g378 (n515, n_9, n514);
  and g379 (n516, \a[3] , \shift[0] );
  and g380 (n517, n_9, n516);
  not g385 (n_212, n519);
  and g386 (n520, n302, n_212);
  and g387 (n521, \a[5] , \shift[0] );
  and g388 (n522, \shift[1] , n521);
  and g389 (n523, \a[6] , n_5);
  and g390 (n524, \shift[1] , n523);
  and g394 (n526, \a[8] , n_5);
  and g395 (n527, n_9, n526);
  and g396 (n528, \a[7] , \shift[0] );
  and g397 (n529, n_9, n528);
  not g402 (n_221, n531);
  and g403 (n532, n315, n_221);
  not g408 (n_224, n534);
  and g409 (n535, n319, n_224);
  and g410 (n536, \a[29] , \shift[0] );
  and g411 (n537, \shift[1] , n536);
  and g412 (n538, \a[30] , n_5);
  and g413 (n539, \shift[1] , n538);
  and g417 (n541, \a[32] , n_5);
  and g418 (n542, n_9, n541);
  and g419 (n543, \a[31] , \shift[0] );
  and g420 (n544, n_9, n543);
  not g425 (n_233, n546);
  and g426 (n547, n275, n_233);
  and g427 (n548, \a[25] , \shift[0] );
  and g428 (n549, \shift[1] , n548);
  and g429 (n550, \a[26] , n_5);
  and g430 (n551, \shift[1] , n550);
  and g434 (n553, \a[28] , n_5);
  and g435 (n554, n_9, n553);
  and g436 (n555, \a[27] , \shift[0] );
  and g437 (n556, n_9, n555);
  not g442 (n_242, n558);
  and g443 (n559, n288, n_242);
  and g447 (n561, \a[17] , \shift[0] );
  and g448 (n562, \shift[1] , n561);
  and g449 (n563, \a[18] , n_5);
  and g450 (n564, \shift[1] , n563);
  and g454 (n566, \a[20] , n_5);
  and g455 (n567, n_9, n566);
  and g456 (n568, \a[19] , \shift[0] );
  and g457 (n569, n_9, n568);
  not g462 (n_253, n571);
  and g463 (n572, n302, n_253);
  and g464 (n573, \a[21] , \shift[0] );
  and g465 (n574, \shift[1] , n573);
  and g466 (n575, \a[22] , n_5);
  and g467 (n576, \shift[1] , n575);
  and g471 (n578, \a[24] , n_5);
  and g472 (n579, n_9, n578);
  and g473 (n580, \a[23] , \shift[0] );
  and g474 (n581, n_9, n580);
  not g479 (n_262, n583);
  and g480 (n584, n315, n_262);
  not g485 (n_265, n586);
  and g486 (n587, n372, n_265);
  and g490 (n589, \a[61] , \shift[0] );
  and g491 (n590, \shift[1] , n589);
  and g492 (n591, \a[62] , n_5);
  and g493 (n592, \shift[1] , n591);
  and g497 (n594, \a[64] , n_5);
  and g498 (n595, n_9, n594);
  and g499 (n596, \a[63] , \shift[0] );
  and g500 (n597, n_9, n596);
  not g505 (n_276, n599);
  and g506 (n600, n275, n_276);
  and g507 (n601, \a[57] , \shift[0] );
  and g508 (n602, \shift[1] , n601);
  and g509 (n603, \a[58] , n_5);
  and g510 (n604, \shift[1] , n603);
  and g514 (n606, \a[60] , n_5);
  and g515 (n607, n_9, n606);
  and g516 (n608, \a[59] , \shift[0] );
  and g517 (n609, n_9, n608);
  not g522 (n_285, n611);
  and g523 (n612, n288, n_285);
  and g527 (n614, \a[49] , \shift[0] );
  and g528 (n615, \shift[1] , n614);
  and g529 (n616, \a[50] , n_5);
  and g530 (n617, \shift[1] , n616);
  and g534 (n619, \a[52] , n_5);
  and g535 (n620, n_9, n619);
  and g536 (n621, \a[51] , \shift[0] );
  and g537 (n622, n_9, n621);
  not g542 (n_296, n624);
  and g543 (n625, n302, n_296);
  and g544 (n626, \a[53] , \shift[0] );
  and g545 (n627, \shift[1] , n626);
  and g546 (n628, \a[54] , n_5);
  and g547 (n629, \shift[1] , n628);
  and g551 (n631, \a[56] , n_5);
  and g552 (n632, n_9, n631);
  and g553 (n633, \a[55] , \shift[0] );
  and g554 (n634, n_9, n633);
  not g559 (n_305, n636);
  and g560 (n637, n315, n_305);
  not g565 (n_308, n639);
  and g566 (n640, n426, n_308);
  and g567 (n641, \a[45] , \shift[0] );
  and g568 (n642, \shift[1] , n641);
  and g569 (n643, \a[46] , n_5);
  and g570 (n644, \shift[1] , n643);
  and g574 (n646, \a[48] , n_5);
  and g575 (n647, n_9, n646);
  and g576 (n648, \a[47] , \shift[0] );
  and g577 (n649, n_9, n648);
  not g582 (n_317, n651);
  and g583 (n652, n275, n_317);
  and g584 (n653, \a[41] , \shift[0] );
  and g585 (n654, \shift[1] , n653);
  and g586 (n655, \a[42] , n_5);
  and g587 (n656, \shift[1] , n655);
  and g591 (n658, \a[44] , n_5);
  and g592 (n659, n_9, n658);
  and g593 (n660, \a[43] , \shift[0] );
  and g594 (n661, n_9, n660);
  not g599 (n_326, n663);
  and g600 (n664, n288, n_326);
  and g604 (n666, \a[33] , \shift[0] );
  and g605 (n667, \shift[1] , n666);
  and g606 (n668, \a[34] , n_5);
  and g607 (n669, \shift[1] , n668);
  and g611 (n671, \a[36] , n_5);
  and g612 (n672, n_9, n671);
  and g613 (n673, \a[35] , \shift[0] );
  and g614 (n674, n_9, n673);
  not g619 (n_337, n676);
  and g620 (n677, n302, n_337);
  and g621 (n678, \a[40] , n_5);
  and g622 (n679, n_9, n678);
  and g623 (n680, \a[37] , \shift[0] );
  and g624 (n681, \shift[1] , n680);
  and g628 (n683, \a[39] , \shift[0] );
  and g629 (n684, n_9, n683);
  and g630 (n685, \a[38] , n_5);
  and g631 (n686, \shift[1] , n685);
  not g636 (n_346, n688);
  and g637 (n689, n315, n_346);
  not g642 (n_349, n691);
  and g643 (n692, n479, n_349);
  not g648 (n_352, n694);
  and g649 (n695, \shift[6] , n_352);
  or g650 (\result[0] , n483, n695);
  and g651 (n697, \a[81] , n_5);
  and g652 (n698, n_9, n697);
  and g653 (n699, \a[78] , \shift[0] );
  and g654 (n700, \shift[1] , n699);
  and g658 (n702, \a[80] , \shift[0] );
  and g659 (n703, n_9, n702);
  and g660 (n704, \a[79] , n_5);
  and g661 (n705, \shift[1] , n704);
  not g666 (n_357, n707);
  and g667 (n708, n275, n_357);
  and g668 (n709, \a[77] , n_5);
  and g669 (n710, n_9, n709);
  and g670 (n711, \a[74] , \shift[0] );
  and g671 (n712, \shift[1] , n711);
  and g675 (n714, \a[76] , \shift[0] );
  and g676 (n715, n_9, n714);
  and g677 (n716, \a[75] , n_5);
  and g678 (n717, \shift[1] , n716);
  not g683 (n_362, n719);
  and g684 (n720, n288, n_362);
  and g688 (n722, \a[69] , n_5);
  and g689 (n723, n_9, n722);
  and g690 (n724, \a[66] , \shift[0] );
  and g691 (n725, \shift[1] , n724);
  and g695 (n727, \a[68] , \shift[0] );
  and g696 (n728, n_9, n727);
  and g697 (n729, \a[67] , n_5);
  and g698 (n730, \shift[1] , n729);
  not g703 (n_369, n732);
  and g704 (n733, n302, n_369);
  and g705 (n734, \a[73] , n_5);
  and g706 (n735, n_9, n734);
  and g707 (n736, \a[70] , \shift[0] );
  and g708 (n737, \shift[1] , n736);
  and g712 (n739, \a[72] , \shift[0] );
  and g713 (n740, n_9, n739);
  and g714 (n741, \a[71] , n_5);
  and g715 (n742, \shift[1] , n741);
  not g720 (n_374, n744);
  and g721 (n745, n315, n_374);
  not g726 (n_377, n747);
  and g727 (n748, n319, n_377);
  and g728 (n749, \a[97] , n_5);
  and g729 (n750, n_9, n749);
  and g730 (n751, \a[94] , \shift[0] );
  and g731 (n752, \shift[1] , n751);
  and g735 (n754, \a[96] , \shift[0] );
  and g736 (n755, n_9, n754);
  and g737 (n756, \a[95] , n_5);
  and g738 (n757, \shift[1] , n756);
  not g743 (n_382, n759);
  and g744 (n760, n275, n_382);
  and g745 (n761, \a[93] , n_5);
  and g746 (n762, n_9, n761);
  and g747 (n763, \a[90] , \shift[0] );
  and g748 (n764, \shift[1] , n763);
  and g752 (n766, \a[92] , \shift[0] );
  and g753 (n767, n_9, n766);
  and g754 (n768, \a[91] , n_5);
  and g755 (n769, \shift[1] , n768);
  not g760 (n_387, n771);
  and g761 (n772, n288, n_387);
  and g765 (n774, \a[85] , n_5);
  and g766 (n775, n_9, n774);
  and g767 (n776, \a[82] , \shift[0] );
  and g768 (n777, \shift[1] , n776);
  and g772 (n779, \a[84] , \shift[0] );
  and g773 (n780, n_9, n779);
  and g774 (n781, \a[83] , n_5);
  and g775 (n782, \shift[1] , n781);
  not g780 (n_394, n784);
  and g781 (n785, n302, n_394);
  and g782 (n786, \a[89] , n_5);
  and g783 (n787, n_9, n786);
  and g784 (n788, \a[86] , \shift[0] );
  and g785 (n789, \shift[1] , n788);
  and g789 (n791, \a[88] , \shift[0] );
  and g790 (n792, n_9, n791);
  and g791 (n793, \a[87] , n_5);
  and g792 (n794, \shift[1] , n793);
  not g797 (n_399, n796);
  and g798 (n797, n315, n_399);
  not g803 (n_402, n799);
  and g804 (n800, n372, n_402);
  and g808 (n802, \a[1] , n_5);
  and g809 (n803, n_9, n802);
  and g810 (n804, \a[126] , \shift[0] );
  and g811 (n805, \shift[1] , n804);
  and g815 (n807, \a[0] , \shift[0] );
  and g816 (n808, n_9, n807);
  and g817 (n809, \a[127] , n_5);
  and g818 (n810, \shift[1] , n809);
  not g823 (n_409, n812);
  and g824 (n813, n275, n_409);
  and g825 (n814, \a[125] , n_5);
  and g826 (n815, n_9, n814);
  and g827 (n816, \a[122] , \shift[0] );
  and g828 (n817, \shift[1] , n816);
  and g832 (n819, \a[124] , \shift[0] );
  and g833 (n820, n_9, n819);
  and g834 (n821, \a[123] , n_5);
  and g835 (n822, \shift[1] , n821);
  not g840 (n_414, n824);
  and g841 (n825, n288, n_414);
  and g845 (n827, \a[117] , n_5);
  and g846 (n828, n_9, n827);
  and g847 (n829, \a[114] , \shift[0] );
  and g848 (n830, \shift[1] , n829);
  and g852 (n832, \a[116] , \shift[0] );
  and g853 (n833, n_9, n832);
  and g854 (n834, \a[115] , n_5);
  and g855 (n835, \shift[1] , n834);
  not g860 (n_421, n837);
  and g861 (n838, n302, n_421);
  and g862 (n839, \a[121] , n_5);
  and g863 (n840, n_9, n839);
  and g864 (n841, \a[118] , \shift[0] );
  and g865 (n842, \shift[1] , n841);
  and g869 (n844, \a[120] , \shift[0] );
  and g870 (n845, n_9, n844);
  and g871 (n846, \a[119] , n_5);
  and g872 (n847, \shift[1] , n846);
  not g877 (n_426, n849);
  and g878 (n850, n315, n_426);
  not g883 (n_429, n852);
  and g884 (n853, n426, n_429);
  and g885 (n854, \a[113] , n_5);
  and g886 (n855, n_9, n854);
  and g887 (n856, \a[110] , \shift[0] );
  and g888 (n857, \shift[1] , n856);
  and g892 (n859, \a[112] , \shift[0] );
  and g893 (n860, n_9, n859);
  and g894 (n861, \a[111] , n_5);
  and g895 (n862, \shift[1] , n861);
  not g900 (n_434, n864);
  and g901 (n865, n275, n_434);
  and g902 (n866, \a[109] , n_5);
  and g903 (n867, n_9, n866);
  and g904 (n868, \a[106] , \shift[0] );
  and g905 (n869, \shift[1] , n868);
  and g909 (n871, \a[108] , \shift[0] );
  and g910 (n872, n_9, n871);
  and g911 (n873, \a[107] , n_5);
  and g912 (n874, \shift[1] , n873);
  not g917 (n_439, n876);
  and g918 (n877, n288, n_439);
  and g922 (n879, \a[101] , n_5);
  and g923 (n880, n_9, n879);
  and g924 (n881, \a[98] , \shift[0] );
  and g925 (n882, \shift[1] , n881);
  and g929 (n884, \a[100] , \shift[0] );
  and g930 (n885, n_9, n884);
  and g931 (n886, \a[99] , n_5);
  and g932 (n887, \shift[1] , n886);
  not g937 (n_446, n889);
  and g938 (n890, n302, n_446);
  and g939 (n891, \a[105] , n_5);
  and g940 (n892, n_9, n891);
  and g941 (n893, \a[102] , \shift[0] );
  and g942 (n894, \shift[1] , n893);
  and g946 (n896, \a[104] , \shift[0] );
  and g947 (n897, n_9, n896);
  and g948 (n898, \a[103] , n_5);
  and g949 (n899, \shift[1] , n898);
  not g954 (n_451, n901);
  and g955 (n902, n315, n_451);
  not g960 (n_454, n904);
  and g961 (n905, n479, n_454);
  not g966 (n_457, n907);
  and g967 (n908, n_182, n_457);
  and g968 (n909, \a[65] , n_5);
  and g969 (n910, n_9, n909);
  and g970 (n911, \a[62] , \shift[0] );
  and g971 (n912, \shift[1] , n911);
  and g975 (n914, \a[64] , \shift[0] );
  and g976 (n915, n_9, n914);
  and g977 (n916, \a[63] , n_5);
  and g978 (n917, \shift[1] , n916);
  not g983 (n_462, n919);
  and g984 (n920, n275, n_462);
  and g985 (n921, \a[61] , n_5);
  and g986 (n922, n_9, n921);
  and g987 (n923, \a[58] , \shift[0] );
  and g988 (n924, \shift[1] , n923);
  and g992 (n926, \a[60] , \shift[0] );
  and g993 (n927, n_9, n926);
  and g994 (n928, \a[59] , n_5);
  and g995 (n929, \shift[1] , n928);
  not g1000 (n_467, n931);
  and g1001 (n932, n288, n_467);
  and g1005 (n934, \a[53] , n_5);
  and g1006 (n935, n_9, n934);
  and g1007 (n936, \a[50] , \shift[0] );
  and g1008 (n937, \shift[1] , n936);
  and g1012 (n939, \a[52] , \shift[0] );
  and g1013 (n940, n_9, n939);
  and g1014 (n941, \a[51] , n_5);
  and g1015 (n942, \shift[1] , n941);
  not g1020 (n_474, n944);
  and g1021 (n945, n302, n_474);
  and g1022 (n946, \a[57] , n_5);
  and g1023 (n947, n_9, n946);
  and g1024 (n948, \a[54] , \shift[0] );
  and g1025 (n949, \shift[1] , n948);
  and g1029 (n951, \a[56] , \shift[0] );
  and g1030 (n952, n_9, n951);
  and g1031 (n953, \a[55] , n_5);
  and g1032 (n954, \shift[1] , n953);
  not g1037 (n_479, n956);
  and g1038 (n957, n315, n_479);
  not g1043 (n_482, n959);
  and g1044 (n960, n426, n_482);
  and g1045 (n961, \a[17] , n_5);
  and g1046 (n962, n_9, n961);
  and g1047 (n963, \a[14] , \shift[0] );
  and g1048 (n964, \shift[1] , n963);
  and g1052 (n966, \a[16] , \shift[0] );
  and g1053 (n967, n_9, n966);
  and g1054 (n968, \a[15] , n_5);
  and g1055 (n969, \shift[1] , n968);
  not g1060 (n_487, n971);
  and g1061 (n972, n275, n_487);
  and g1062 (n973, \a[13] , n_5);
  and g1063 (n974, n_9, n973);
  and g1064 (n975, \a[10] , \shift[0] );
  and g1065 (n976, \shift[1] , n975);
  and g1069 (n978, \a[12] , \shift[0] );
  and g1070 (n979, n_9, n978);
  and g1071 (n980, \a[11] , n_5);
  and g1072 (n981, \shift[1] , n980);
  not g1077 (n_492, n983);
  and g1078 (n984, n288, n_492);
  and g1082 (n986, \a[5] , n_5);
  and g1083 (n987, n_9, n986);
  and g1084 (n988, \a[2] , \shift[0] );
  and g1085 (n989, \shift[1] , n988);
  and g1089 (n991, \a[4] , \shift[0] );
  and g1090 (n992, n_9, n991);
  and g1091 (n993, \a[3] , n_5);
  and g1092 (n994, \shift[1] , n993);
  not g1097 (n_499, n996);
  and g1098 (n997, n302, n_499);
  and g1099 (n998, \a[9] , n_5);
  and g1100 (n999, n_9, n998);
  and g1101 (n1000, \a[6] , \shift[0] );
  and g1102 (n1001, \shift[1] , n1000);
  and g1106 (n1003, \a[8] , \shift[0] );
  and g1107 (n1004, n_9, n1003);
  and g1108 (n1005, \a[7] , n_5);
  and g1109 (n1006, \shift[1] , n1005);
  not g1114 (n_504, n1008);
  and g1115 (n1009, n315, n_504);
  not g1120 (n_507, n1011);
  and g1121 (n1012, n319, n_507);
  and g1125 (n1014, \a[49] , n_5);
  and g1126 (n1015, n_9, n1014);
  and g1127 (n1016, \a[46] , \shift[0] );
  and g1128 (n1017, \shift[1] , n1016);
  and g1132 (n1019, \a[48] , \shift[0] );
  and g1133 (n1020, n_9, n1019);
  and g1134 (n1021, \a[47] , n_5);
  and g1135 (n1022, \shift[1] , n1021);
  not g1140 (n_514, n1024);
  and g1141 (n1025, n275, n_514);
  and g1142 (n1026, \a[42] , \shift[0] );
  and g1143 (n1027, \shift[1] , n1026);
  and g1144 (n1028, \a[43] , n_5);
  and g1145 (n1029, \shift[1] , n1028);
  and g1149 (n1031, \a[45] , n_5);
  and g1150 (n1032, n_9, n1031);
  and g1151 (n1033, \a[44] , \shift[0] );
  and g1152 (n1034, n_9, n1033);
  not g1157 (n_519, n1036);
  and g1158 (n1037, n288, n_519);
  and g1162 (n1039, \a[37] , n_5);
  and g1163 (n1040, n_9, n1039);
  and g1164 (n1041, \a[34] , \shift[0] );
  and g1165 (n1042, \shift[1] , n1041);
  and g1169 (n1044, \a[36] , \shift[0] );
  and g1170 (n1045, n_9, n1044);
  and g1171 (n1046, \a[35] , n_5);
  and g1172 (n1047, \shift[1] , n1046);
  not g1177 (n_526, n1049);
  and g1178 (n1050, n302, n_526);
  and g1179 (n1051, \a[41] , n_5);
  and g1180 (n1052, n_9, n1051);
  and g1181 (n1053, \a[40] , \shift[0] );
  and g1182 (n1054, n_9, n1053);
  and g1186 (n1056, \a[39] , n_5);
  and g1187 (n1057, \shift[1] , n1056);
  and g1188 (n1058, \a[38] , \shift[0] );
  and g1189 (n1059, \shift[1] , n1058);
  not g1194 (n_531, n1061);
  and g1195 (n1062, n315, n_531);
  not g1200 (n_534, n1064);
  and g1201 (n1065, n479, n_534);
  and g1202 (n1066, \a[33] , n_5);
  and g1203 (n1067, n_9, n1066);
  and g1204 (n1068, \a[30] , \shift[0] );
  and g1205 (n1069, \shift[1] , n1068);
  and g1209 (n1071, \a[32] , \shift[0] );
  and g1210 (n1072, n_9, n1071);
  and g1211 (n1073, \a[31] , n_5);
  and g1212 (n1074, \shift[1] , n1073);
  not g1217 (n_539, n1076);
  and g1218 (n1077, n275, n_539);
  and g1219 (n1078, \a[29] , n_5);
  and g1220 (n1079, n_9, n1078);
  and g1221 (n1080, \a[26] , \shift[0] );
  and g1222 (n1081, \shift[1] , n1080);
  and g1226 (n1083, \a[28] , \shift[0] );
  and g1227 (n1084, n_9, n1083);
  and g1228 (n1085, \a[27] , n_5);
  and g1229 (n1086, \shift[1] , n1085);
  not g1234 (n_544, n1088);
  and g1235 (n1089, n288, n_544);
  and g1239 (n1091, \a[21] , n_5);
  and g1240 (n1092, n_9, n1091);
  and g1241 (n1093, \a[18] , \shift[0] );
  and g1242 (n1094, \shift[1] , n1093);
  and g1246 (n1096, \a[20] , \shift[0] );
  and g1247 (n1097, n_9, n1096);
  and g1248 (n1098, \a[19] , n_5);
  and g1249 (n1099, \shift[1] , n1098);
  not g1254 (n_551, n1101);
  and g1255 (n1102, n302, n_551);
  and g1256 (n1103, \a[25] , n_5);
  and g1257 (n1104, n_9, n1103);
  and g1258 (n1105, \a[22] , \shift[0] );
  and g1259 (n1106, \shift[1] , n1105);
  and g1263 (n1108, \a[24] , \shift[0] );
  and g1264 (n1109, n_9, n1108);
  and g1265 (n1110, \a[23] , n_5);
  and g1266 (n1111, \shift[1] , n1110);
  not g1271 (n_556, n1113);
  and g1272 (n1114, n315, n_556);
  not g1277 (n_559, n1116);
  and g1278 (n1117, n372, n_559);
  not g1283 (n_562, n1119);
  and g1284 (n1120, \shift[6] , n_562);
  or g1285 (\result[1] , n908, n1120);
  and g1286 (n1122, n_9, n346);
  and g1287 (n1123, n_9, n348);
  and g1291 (n1125, \shift[1] , n269);
  and g1292 (n1126, \shift[1] , n271);
  not g1297 (n_567, n1128);
  and g1298 (n1129, n275, n_567);
  and g1299 (n1130, n_9, n264);
  and g1300 (n1131, n_9, n266);
  and g1304 (n1133, \shift[1] , n282);
  and g1305 (n1134, \shift[1] , n284);
  not g1310 (n_572, n1136);
  and g1311 (n1137, n288, n_572);
  and g1315 (n1139, n_9, n304);
  and g1316 (n1140, n_9, n306);
  and g1320 (n1142, \shift[1] , n296);
  and g1321 (n1143, \shift[1] , n298);
  not g1326 (n_579, n1145);
  and g1327 (n1146, n302, n_579);
  and g1328 (n1147, n_9, n277);
  and g1329 (n1148, n_9, n279);
  and g1333 (n1150, \shift[1] , n309);
  and g1334 (n1151, \shift[1] , n311);
  not g1339 (n_584, n1153);
  and g1340 (n1154, n315, n_584);
  not g1345 (n_587, n1156);
  and g1346 (n1157, n319, n_587);
  and g1347 (n1158, n_9, n453);
  and g1348 (n1159, n_9, n455);
  and g1352 (n1161, \shift[1] , n326);
  and g1353 (n1162, \shift[1] , n328);
  not g1358 (n_592, n1164);
  and g1359 (n1165, n275, n_592);
  and g1360 (n1166, n_9, n321);
  and g1361 (n1167, n_9, n323);
  and g1365 (n1169, \shift[1] , n338);
  and g1366 (n1170, \shift[1] , n340);
  not g1371 (n_597, n1172);
  and g1372 (n1173, n288, n_597);
  and g1376 (n1175, n_9, n358);
  and g1377 (n1176, n_9, n360);
  and g1381 (n1178, \shift[1] , n351);
  and g1382 (n1179, \shift[1] , n353);
  not g1387 (n_604, n1181);
  and g1388 (n1182, n302, n_604);
  and g1389 (n1183, n_9, n333);
  and g1390 (n1184, n_9, n335);
  and g1394 (n1186, \shift[1] , n363);
  and g1395 (n1187, \shift[1] , n365);
  not g1400 (n_609, n1189);
  and g1401 (n1190, n315, n_609);
  not g1406 (n_612, n1192);
  and g1407 (n1193, n372, n_612);
  and g1411 (n1195, n_9, n509);
  and g1412 (n1196, n_9, n511);
  and g1416 (n1198, \shift[1] , n380);
  and g1417 (n1199, \shift[1] , n382);
  not g1422 (n_619, n1201);
  and g1423 (n1202, n275, n_619);
  and g1424 (n1203, n_9, n375);
  and g1425 (n1204, n_9, n377);
  and g1429 (n1206, \shift[1] , n392);
  and g1430 (n1207, \shift[1] , n394);
  not g1435 (n_624, n1209);
  and g1436 (n1210, n288, n_624);
  and g1440 (n1212, n_9, n412);
  and g1441 (n1213, n_9, n414);
  and g1445 (n1215, \shift[1] , n405);
  and g1446 (n1216, \shift[1] , n407);
  not g1451 (n_631, n1218);
  and g1452 (n1219, n302, n_631);
  and g1453 (n1220, n_9, n387);
  and g1454 (n1221, n_9, n389);
  and g1458 (n1223, \shift[1] , n417);
  and g1459 (n1224, \shift[1] , n419);
  not g1464 (n_636, n1226);
  and g1465 (n1227, n315, n_636);
  not g1470 (n_639, n1229);
  and g1471 (n1230, n426, n_639);
  and g1472 (n1231, n_9, n400);
  and g1473 (n1232, n_9, n402);
  and g1477 (n1234, \shift[1] , n433);
  and g1478 (n1235, \shift[1] , n435);
  not g1483 (n_644, n1237);
  and g1484 (n1238, n275, n_644);
  and g1485 (n1239, n_9, n428);
  and g1486 (n1240, n_9, n430);
  and g1490 (n1242, \shift[1] , n445);
  and g1491 (n1243, \shift[1] , n447);
  not g1496 (n_649, n1245);
  and g1497 (n1246, n288, n_649);
  and g1501 (n1248, n_9, n465);
  and g1502 (n1249, n_9, n467);
  and g1506 (n1251, \shift[1] , n458);
  and g1507 (n1252, \shift[1] , n460);
  not g1512 (n_656, n1254);
  and g1513 (n1255, n302, n_656);
  and g1514 (n1256, n_9, n440);
  and g1515 (n1257, n_9, n442);
  and g1519 (n1259, \shift[1] , n470);
  and g1520 (n1260, \shift[1] , n472);
  not g1525 (n_661, n1262);
  and g1526 (n1263, n315, n_661);
  not g1531 (n_664, n1265);
  and g1532 (n1266, n479, n_664);
  not g1537 (n_667, n1268);
  and g1538 (n1269, n_182, n_667);
  and g1539 (n1270, n_9, n291);
  and g1540 (n1271, n_9, n293);
  and g1544 (n1273, \shift[1] , n594);
  and g1545 (n1274, \shift[1] , n596);
  not g1550 (n_672, n1276);
  and g1551 (n1277, n275, n_672);
  and g1552 (n1278, n_9, n589);
  and g1553 (n1279, n_9, n591);
  and g1557 (n1281, \shift[1] , n606);
  and g1558 (n1282, \shift[1] , n608);
  not g1563 (n_677, n1284);
  and g1564 (n1285, n288, n_677);
  and g1568 (n1287, n_9, n626);
  and g1569 (n1288, n_9, n628);
  and g1573 (n1290, \shift[1] , n619);
  and g1574 (n1291, \shift[1] , n621);
  not g1579 (n_684, n1293);
  and g1580 (n1294, n302, n_684);
  and g1581 (n1295, n_9, n601);
  and g1582 (n1296, n_9, n603);
  and g1586 (n1298, \shift[1] , n631);
  and g1587 (n1299, \shift[1] , n633);
  not g1592 (n_689, n1301);
  and g1593 (n1302, n315, n_689);
  not g1598 (n_692, n1304);
  and g1599 (n1305, n426, n_692);
  and g1600 (n1306, n_9, n561);
  and g1601 (n1307, n_9, n563);
  and g1605 (n1309, \shift[1] , n489);
  and g1606 (n1310, \shift[1] , n491);
  not g1611 (n_697, n1312);
  and g1612 (n1313, n275, n_697);
  and g1613 (n1314, n_9, n484);
  and g1614 (n1315, n_9, n486);
  and g1618 (n1317, \shift[1] , n501);
  and g1619 (n1318, \shift[1] , n503);
  not g1624 (n_702, n1320);
  and g1625 (n1321, n288, n_702);
  and g1629 (n1323, n_9, n521);
  and g1630 (n1324, n_9, n523);
  and g1634 (n1326, \shift[1] , n514);
  and g1635 (n1327, \shift[1] , n516);
  not g1640 (n_709, n1329);
  and g1641 (n1330, n302, n_709);
  and g1642 (n1331, n_9, n496);
  and g1643 (n1332, n_9, n498);
  and g1647 (n1334, \shift[1] , n526);
  and g1648 (n1335, \shift[1] , n528);
  not g1653 (n_714, n1337);
  and g1654 (n1338, n315, n_714);
  not g1659 (n_717, n1340);
  and g1660 (n1341, n319, n_717);
  and g1664 (n1343, n_9, n614);
  and g1665 (n1344, n_9, n616);
  and g1669 (n1346, \shift[1] , n646);
  and g1670 (n1347, \shift[1] , n648);
  not g1675 (n_724, n1349);
  and g1676 (n1350, n275, n_724);
  and g1677 (n1351, \shift[1] , n660);
  and g1678 (n1352, \shift[1] , n658);
  and g1682 (n1354, n_9, n643);
  and g1683 (n1355, n_9, n641);
  not g1688 (n_729, n1357);
  and g1689 (n1358, n288, n_729);
  and g1693 (n1360, n_9, n680);
  and g1694 (n1361, n_9, n685);
  and g1698 (n1363, \shift[1] , n671);
  and g1699 (n1364, \shift[1] , n673);
  not g1704 (n_736, n1366);
  and g1705 (n1367, n302, n_736);
  and g1706 (n1368, n_9, n653);
  and g1707 (n1369, n_9, n655);
  and g1711 (n1371, \shift[1] , n683);
  and g1712 (n1372, \shift[1] , n678);
  not g1717 (n_741, n1374);
  and g1718 (n1375, n315, n_741);
  not g1723 (n_744, n1377);
  and g1724 (n1378, n479, n_744);
  and g1725 (n1379, n_9, n666);
  and g1726 (n1380, n_9, n668);
  and g1730 (n1382, \shift[1] , n541);
  and g1731 (n1383, \shift[1] , n543);
  not g1736 (n_749, n1385);
  and g1737 (n1386, n275, n_749);
  and g1738 (n1387, n_9, n536);
  and g1739 (n1388, n_9, n538);
  and g1743 (n1390, \shift[1] , n553);
  and g1744 (n1391, \shift[1] , n555);
  not g1749 (n_754, n1393);
  and g1750 (n1394, n288, n_754);
  and g1754 (n1396, n_9, n573);
  and g1755 (n1397, n_9, n575);
  and g1759 (n1399, \shift[1] , n566);
  and g1760 (n1400, \shift[1] , n568);
  not g1765 (n_761, n1402);
  and g1766 (n1403, n302, n_761);
  and g1767 (n1404, n_9, n548);
  and g1768 (n1405, n_9, n550);
  and g1772 (n1407, \shift[1] , n578);
  and g1773 (n1408, \shift[1] , n580);
  not g1778 (n_766, n1410);
  and g1779 (n1411, n315, n_766);
  not g1784 (n_769, n1413);
  and g1785 (n1414, n372, n_769);
  not g1790 (n_772, n1416);
  and g1791 (n1417, \shift[6] , n_772);
  or g1792 (\result[2] , n1269, n1417);
  and g1793 (n1419, \shift[1] , n854);
  and g1794 (n1420, n_9, n829);
  and g1798 (n1422, \shift[1] , n859);
  and g1799 (n1423, n_9, n834);
  not g1804 (n_777, n1425);
  and g1805 (n1426, n275, n_777);
  and g1806 (n1427, \shift[1] , n866);
  and g1807 (n1428, n_9, n856);
  and g1811 (n1430, \shift[1] , n871);
  and g1812 (n1431, n_9, n861);
  not g1817 (n_782, n1433);
  and g1818 (n1434, n288, n_782);
  and g1822 (n1436, \shift[1] , n879);
  and g1823 (n1437, n_9, n893);
  and g1827 (n1439, \shift[1] , n884);
  and g1828 (n1440, n_9, n898);
  not g1833 (n_789, n1442);
  and g1834 (n1443, n302, n_789);
  and g1835 (n1444, \shift[1] , n891);
  and g1836 (n1445, n_9, n868);
  and g1840 (n1447, \shift[1] , n896);
  and g1841 (n1448, n_9, n873);
  not g1846 (n_794, n1450);
  and g1847 (n1451, n315, n_794);
  not g1852 (n_797, n1453);
  and g1853 (n1454, n479, n_797);
  and g1854 (n1455, \shift[1] , n749);
  and g1855 (n1456, n_9, n881);
  and g1859 (n1458, \shift[1] , n754);
  and g1860 (n1459, n_9, n886);
  not g1865 (n_802, n1461);
  and g1866 (n1462, n275, n_802);
  and g1867 (n1463, \shift[1] , n761);
  and g1868 (n1464, n_9, n751);
  and g1872 (n1466, \shift[1] , n766);
  and g1873 (n1467, n_9, n756);
  not g1878 (n_807, n1469);
  and g1879 (n1470, n288, n_807);
  and g1883 (n1472, \shift[1] , n774);
  and g1884 (n1473, n_9, n788);
  and g1888 (n1475, \shift[1] , n779);
  and g1889 (n1476, n_9, n793);
  not g1894 (n_814, n1478);
  and g1895 (n1479, n302, n_814);
  and g1896 (n1480, \shift[1] , n786);
  and g1897 (n1481, n_9, n763);
  and g1901 (n1483, \shift[1] , n791);
  and g1902 (n1484, n_9, n768);
  not g1907 (n_819, n1486);
  and g1908 (n1487, n315, n_819);
  not g1913 (n_822, n1489);
  and g1914 (n1490, n372, n_822);
  and g1918 (n1492, \shift[1] , n802);
  and g1919 (n1493, n_9, n988);
  and g1923 (n1495, \shift[1] , n807);
  and g1924 (n1496, n_9, n993);
  not g1929 (n_829, n1498);
  and g1930 (n1499, n275, n_829);
  and g1931 (n1500, \shift[1] , n814);
  and g1932 (n1501, n_9, n804);
  and g1936 (n1503, \shift[1] , n819);
  and g1937 (n1504, n_9, n809);
  not g1942 (n_834, n1506);
  and g1943 (n1507, n288, n_834);
  and g1947 (n1509, \shift[1] , n827);
  and g1948 (n1510, n_9, n841);
  and g1952 (n1512, \shift[1] , n832);
  and g1953 (n1513, n_9, n846);
  not g1958 (n_841, n1515);
  and g1959 (n1516, n302, n_841);
  and g1960 (n1517, \shift[1] , n839);
  and g1961 (n1518, n_9, n816);
  and g1965 (n1520, \shift[1] , n844);
  and g1966 (n1521, n_9, n821);
  not g1971 (n_846, n1523);
  and g1972 (n1524, n315, n_846);
  not g1977 (n_849, n1526);
  and g1978 (n1527, n426, n_849);
  and g1979 (n1528, \shift[1] , n697);
  and g1980 (n1529, n_9, n776);
  and g1984 (n1531, \shift[1] , n702);
  and g1985 (n1532, n_9, n781);
  not g1990 (n_854, n1534);
  and g1991 (n1535, n275, n_854);
  and g1992 (n1536, \shift[1] , n709);
  and g1993 (n1537, n_9, n699);
  and g1997 (n1539, \shift[1] , n714);
  and g1998 (n1540, n_9, n704);
  not g2003 (n_859, n1542);
  and g2004 (n1543, n288, n_859);
  and g2008 (n1545, \shift[1] , n722);
  and g2009 (n1546, n_9, n736);
  and g2013 (n1548, \shift[1] , n727);
  and g2014 (n1549, n_9, n741);
  not g2019 (n_866, n1551);
  and g2020 (n1552, n302, n_866);
  and g2021 (n1553, \shift[1] , n734);
  and g2022 (n1554, n_9, n711);
  and g2026 (n1556, \shift[1] , n739);
  and g2027 (n1557, n_9, n716);
  not g2032 (n_871, n1559);
  and g2033 (n1560, n315, n_871);
  not g2038 (n_874, n1562);
  and g2039 (n1563, n319, n_874);
  not g2044 (n_877, n1565);
  and g2045 (n1566, n_182, n_877);
  and g2046 (n1567, \shift[1] , n909);
  and g2047 (n1568, n_9, n724);
  and g2051 (n1570, \shift[1] , n914);
  and g2052 (n1571, n_9, n729);
  not g2057 (n_882, n1573);
  and g2058 (n1574, n275, n_882);
  and g2059 (n1575, \shift[1] , n921);
  and g2060 (n1576, n_9, n911);
  and g2064 (n1578, \shift[1] , n926);
  and g2065 (n1579, n_9, n916);
  not g2070 (n_887, n1581);
  and g2071 (n1582, n288, n_887);
  and g2075 (n1584, \shift[1] , n934);
  and g2076 (n1585, n_9, n948);
  and g2080 (n1587, \shift[1] , n939);
  and g2081 (n1588, n_9, n953);
  not g2086 (n_894, n1590);
  and g2087 (n1591, n302, n_894);
  and g2088 (n1592, \shift[1] , n946);
  and g2089 (n1593, n_9, n923);
  and g2093 (n1595, \shift[1] , n951);
  and g2094 (n1596, n_9, n928);
  not g2099 (n_899, n1598);
  and g2100 (n1599, n315, n_899);
  not g2105 (n_902, n1601);
  and g2106 (n1602, n426, n_902);
  and g2107 (n1603, \shift[1] , n1014);
  and g2108 (n1604, n_9, n936);
  and g2112 (n1606, \shift[1] , n1019);
  and g2113 (n1607, n_9, n941);
  not g2118 (n_907, n1609);
  and g2119 (n1610, n275, n_907);
  and g2120 (n1611, \shift[1] , n1033);
  and g2121 (n1612, \shift[1] , n1031);
  and g2125 (n1614, n_9, n1021);
  and g2126 (n1615, n_9, n1016);
  not g2131 (n_912, n1617);
  and g2132 (n1618, n288, n_912);
  and g2136 (n1620, \shift[1] , n1039);
  and g2137 (n1621, n_9, n1058);
  and g2141 (n1623, \shift[1] , n1044);
  and g2142 (n1624, n_9, n1056);
  not g2147 (n_919, n1626);
  and g2148 (n1627, n302, n_919);
  and g2149 (n1628, \shift[1] , n1051);
  and g2150 (n1629, n_9, n1026);
  and g2154 (n1631, \shift[1] , n1053);
  and g2155 (n1632, n_9, n1028);
  not g2160 (n_924, n1634);
  and g2161 (n1635, n315, n_924);
  not g2166 (n_927, n1637);
  and g2167 (n1638, n479, n_927);
  and g2171 (n1640, \shift[1] , n961);
  and g2172 (n1641, n_9, n1093);
  and g2176 (n1643, \shift[1] , n966);
  and g2177 (n1644, n_9, n1098);
  not g2182 (n_934, n1646);
  and g2183 (n1647, n275, n_934);
  and g2184 (n1648, \shift[1] , n973);
  and g2185 (n1649, n_9, n963);
  and g2189 (n1651, \shift[1] , n978);
  and g2190 (n1652, n_9, n968);
  not g2195 (n_939, n1654);
  and g2196 (n1655, n288, n_939);
  and g2200 (n1657, \shift[1] , n986);
  and g2201 (n1658, n_9, n1000);
  and g2205 (n1660, \shift[1] , n991);
  and g2206 (n1661, n_9, n1005);
  not g2211 (n_946, n1663);
  and g2212 (n1664, n302, n_946);
  and g2213 (n1665, \shift[1] , n998);
  and g2214 (n1666, n_9, n975);
  and g2218 (n1668, \shift[1] , n1003);
  and g2219 (n1669, n_9, n980);
  not g2224 (n_951, n1671);
  and g2225 (n1672, n315, n_951);
  not g2230 (n_954, n1674);
  and g2231 (n1675, n319, n_954);
  and g2232 (n1676, \shift[1] , n1066);
  and g2233 (n1677, n_9, n1041);
  and g2237 (n1679, \shift[1] , n1071);
  and g2238 (n1680, n_9, n1046);
  not g2243 (n_959, n1682);
  and g2244 (n1683, n275, n_959);
  and g2245 (n1684, \shift[1] , n1078);
  and g2246 (n1685, n_9, n1068);
  and g2250 (n1687, \shift[1] , n1083);
  and g2251 (n1688, n_9, n1073);
  not g2256 (n_964, n1690);
  and g2257 (n1691, n288, n_964);
  and g2261 (n1693, \shift[1] , n1091);
  and g2262 (n1694, n_9, n1105);
  and g2266 (n1696, \shift[1] , n1096);
  and g2267 (n1697, n_9, n1110);
  not g2272 (n_971, n1699);
  and g2273 (n1700, n302, n_971);
  and g2274 (n1701, \shift[1] , n1103);
  and g2275 (n1702, n_9, n1080);
  and g2279 (n1704, \shift[1] , n1108);
  and g2280 (n1705, n_9, n1085);
  not g2285 (n_976, n1707);
  and g2286 (n1708, n315, n_976);
  not g2291 (n_979, n1710);
  and g2292 (n1711, n372, n_979);
  not g2297 (n_982, n1713);
  and g2298 (n1714, \shift[6] , n_982);
  or g2299 (\result[3] , n1566, n1714);
  and g2300 (n1716, n275, n_80);
  and g2301 (n1717, n_17, n288);
  and g2305 (n1719, n302, n_46);
  and g2306 (n1720, n_26, n315);
  not g2311 (n_987, n1722);
  and g2312 (n1723, n319, n_987);
  and g2313 (n1724, n275, n_166);
  and g2314 (n1725, n288, n_60);
  and g2318 (n1727, n302, n_89);
  and g2319 (n1728, n315, n_69);
  not g2324 (n_992, n1730);
  and g2325 (n1731, n372, n_992);
  and g2329 (n1733, n275, n_212);
  and g2330 (n1734, n288, n_104);
  and g2334 (n1736, n302, n_133);
  and g2335 (n1737, n315, n_113);
  not g2340 (n_999, n1739);
  and g2341 (n1740, n426, n_999);
  and g2342 (n1741, n275, n_124);
  and g2343 (n1742, n288, n_146);
  and g2347 (n1744, n302, n_175);
  and g2348 (n1745, n315, n_155);
  not g2353 (n_1004, n1747);
  and g2354 (n1748, n479, n_1004);
  not g2359 (n_1007, n1750);
  and g2360 (n1751, n_182, n_1007);
  and g2361 (n1752, n275, n_296);
  and g2362 (n1753, n288, n_317);
  and g2366 (n1755, n302, n_346);
  and g2367 (n1756, n315, n_326);
  not g2372 (n_1012, n1758);
  and g2373 (n1759, n479, n_1012);
  and g2374 (n1760, n275, n_37);
  and g2375 (n1761, n288, n_276);
  and g2379 (n1763, n302, n_305);
  and g2380 (n1764, n315, n_285);
  not g2385 (n_1017, n1766);
  and g2386 (n1767, n426, n_1017);
  and g2390 (n1769, n275, n_337);
  and g2391 (n1770, n288, n_233);
  and g2395 (n1772, n302, n_262);
  and g2396 (n1773, n315, n_242);
  not g2401 (n_1024, n1775);
  and g2402 (n1776, n372, n_1024);
  and g2403 (n1777, n275, n_253);
  and g2404 (n1778, n288, n_192);
  and g2408 (n1780, n302, n_221);
  and g2409 (n1781, n315, n_201);
  not g2414 (n_1029, n1783);
  and g2415 (n1784, n319, n_1029);
  not g2420 (n_1032, n1786);
  and g2421 (n1787, \shift[6] , n_1032);
  or g2422 (\result[4] , n1751, n1787);
  and g2423 (n1789, n275, n_394);
  and g2424 (n1790, n288, n_357);
  and g2428 (n1792, n302, n_374);
  and g2429 (n1793, n315, n_362);
  not g2434 (n_1037, n1795);
  and g2435 (n1796, n319, n_1037);
  and g2436 (n1797, n275, n_446);
  and g2437 (n1798, n288, n_382);
  and g2441 (n1800, n302, n_399);
  and g2442 (n1801, n315, n_387);
  not g2447 (n_1042, n1803);
  and g2448 (n1804, n372, n_1042);
  and g2452 (n1806, n275, n_499);
  and g2453 (n1807, n288, n_409);
  and g2457 (n1809, n302, n_426);
  and g2458 (n1810, n315, n_414);
  not g2463 (n_1049, n1812);
  and g2464 (n1813, n426, n_1049);
  and g2465 (n1814, n275, n_421);
  and g2466 (n1815, n288, n_434);
  and g2470 (n1817, n302, n_451);
  and g2471 (n1818, n315, n_439);
  not g2476 (n_1054, n1820);
  and g2477 (n1821, n479, n_1054);
  not g2482 (n_1057, n1823);
  and g2483 (n1824, n_182, n_1057);
  and g2484 (n1825, n275, n_474);
  and g2485 (n1826, n288, n_514);
  and g2489 (n1828, n302, n_531);
  and g2490 (n1829, n315, n_519);
  not g2495 (n_1062, n1831);
  and g2496 (n1832, n479, n_1062);
  and g2497 (n1833, n275, n_369);
  and g2498 (n1834, n288, n_462);
  and g2502 (n1836, n302, n_479);
  and g2503 (n1837, n315, n_467);
  not g2508 (n_1067, n1839);
  and g2509 (n1840, n426, n_1067);
  and g2513 (n1842, n275, n_526);
  and g2514 (n1843, n288, n_539);
  and g2518 (n1845, n302, n_556);
  and g2519 (n1846, n315, n_544);
  not g2524 (n_1074, n1848);
  and g2525 (n1849, n372, n_1074);
  and g2526 (n1850, n275, n_551);
  and g2527 (n1851, n288, n_487);
  and g2531 (n1853, n302, n_504);
  and g2532 (n1854, n315, n_492);
  not g2537 (n_1079, n1856);
  and g2538 (n1857, n319, n_1079);
  not g2543 (n_1082, n1859);
  and g2544 (n1860, \shift[6] , n_1082);
  or g2545 (\result[5] , n1824, n1860);
  and g2546 (n1862, n275, n_604);
  and g2547 (n1863, n288, n_567);
  and g2551 (n1865, n302, n_584);
  and g2552 (n1866, n315, n_572);
  not g2557 (n_1087, n1868);
  and g2558 (n1869, n319, n_1087);
  and g2559 (n1870, n275, n_656);
  and g2560 (n1871, n288, n_592);
  and g2564 (n1873, n302, n_609);
  and g2565 (n1874, n315, n_597);
  not g2570 (n_1092, n1876);
  and g2571 (n1877, n372, n_1092);
  and g2575 (n1879, n275, n_709);
  and g2576 (n1880, n288, n_619);
  and g2580 (n1882, n302, n_636);
  and g2581 (n1883, n315, n_624);
  not g2586 (n_1099, n1885);
  and g2587 (n1886, n426, n_1099);
  and g2588 (n1887, n275, n_631);
  and g2589 (n1888, n288, n_644);
  and g2593 (n1890, n302, n_661);
  and g2594 (n1891, n315, n_649);
  not g2599 (n_1104, n1893);
  and g2600 (n1894, n479, n_1104);
  not g2605 (n_1107, n1896);
  and g2606 (n1897, n_182, n_1107);
  and g2607 (n1898, n275, n_684);
  and g2608 (n1899, n288, n_724);
  and g2612 (n1901, n302, n_741);
  and g2613 (n1902, n315, n_729);
  not g2618 (n_1112, n1904);
  and g2619 (n1905, n479, n_1112);
  and g2620 (n1906, n275, n_579);
  and g2621 (n1907, n288, n_672);
  and g2625 (n1909, n302, n_689);
  and g2626 (n1910, n315, n_677);
  not g2631 (n_1117, n1912);
  and g2632 (n1913, n426, n_1117);
  and g2636 (n1915, n275, n_736);
  and g2637 (n1916, n288, n_749);
  and g2641 (n1918, n302, n_766);
  and g2642 (n1919, n315, n_754);
  not g2647 (n_1124, n1921);
  and g2648 (n1922, n372, n_1124);
  and g2649 (n1923, n275, n_761);
  and g2650 (n1924, n288, n_697);
  and g2654 (n1926, n302, n_714);
  and g2655 (n1927, n315, n_702);
  not g2660 (n_1129, n1929);
  and g2661 (n1930, n319, n_1129);
  not g2666 (n_1132, n1932);
  and g2667 (n1933, \shift[6] , n_1132);
  or g2668 (\result[6] , n1897, n1933);
  and g2669 (n1935, n275, n_814);
  and g2670 (n1936, n288, n_854);
  and g2674 (n1938, n302, n_871);
  and g2675 (n1939, n315, n_859);
  not g2680 (n_1137, n1941);
  and g2681 (n1942, n319, n_1137);
  and g2682 (n1943, n275, n_789);
  and g2683 (n1944, n288, n_802);
  and g2687 (n1946, n302, n_819);
  and g2688 (n1947, n315, n_807);
  not g2693 (n_1142, n1949);
  and g2694 (n1950, n372, n_1142);
  and g2698 (n1952, n275, n_946);
  and g2699 (n1953, n288, n_829);
  and g2703 (n1955, n302, n_846);
  and g2704 (n1956, n315, n_834);
  not g2709 (n_1149, n1958);
  and g2710 (n1959, n426, n_1149);
  and g2711 (n1960, n275, n_841);
  and g2712 (n1961, n288, n_777);
  and g2716 (n1963, n302, n_794);
  and g2717 (n1964, n315, n_782);
  not g2722 (n_1154, n1966);
  and g2723 (n1967, n479, n_1154);
  not g2728 (n_1157, n1969);
  and g2729 (n1970, n_182, n_1157);
  and g2730 (n1971, n288, n_907);
  and g2731 (n1972, n315, n_912);
  and g2735 (n1974, n302, n_924);
  and g2736 (n1975, n275, n_894);
  not g2741 (n_1162, n1977);
  and g2742 (n1978, n479, n_1162);
  and g2743 (n1979, n275, n_866);
  and g2744 (n1980, n288, n_882);
  and g2748 (n1982, n302, n_899);
  and g2749 (n1983, n315, n_887);
  not g2754 (n_1167, n1985);
  and g2755 (n1986, n426, n_1167);
  and g2759 (n1988, n275, n_919);
  and g2760 (n1989, n288, n_959);
  and g2764 (n1991, n302, n_976);
  and g2765 (n1992, n315, n_964);
  not g2770 (n_1174, n1994);
  and g2771 (n1995, n372, n_1174);
  and g2772 (n1996, n275, n_971);
  and g2773 (n1997, n288, n_934);
  and g2777 (n1999, n302, n_951);
  and g2778 (n2000, n315, n_939);
  not g2783 (n_1179, n2002);
  and g2784 (n2003, n319, n_1179);
  not g2789 (n_1182, n2005);
  and g2790 (n2006, \shift[6] , n_1182);
  or g2791 (\result[7] , n1970, n2006);
  and g2792 (n2008, n275, n_89);
  and g2793 (n2009, n288, n_80);
  and g2797 (n2011, n_26, n302);
  and g2798 (n2012, n_17, n315);
  not g2803 (n_1187, n2014);
  and g2804 (n2015, n319, n_1187);
  and g2805 (n2016, n275, n_175);
  and g2806 (n2017, n288, n_166);
  and g2810 (n2019, n302, n_69);
  and g2811 (n2020, n315, n_60);
  not g2816 (n_1192, n2022);
  and g2817 (n2023, n372, n_1192);
  and g2821 (n2025, n275, n_221);
  and g2822 (n2026, n288, n_212);
  and g2826 (n2028, n302, n_113);
  and g2827 (n2029, n315, n_104);
  not g2832 (n_1199, n2031);
  and g2833 (n2032, n426, n_1199);
  and g2834 (n2033, n275, n_133);
  and g2835 (n2034, n288, n_124);
  and g2839 (n2036, n302, n_155);
  and g2840 (n2037, n315, n_146);
  not g2845 (n_1204, n2039);
  and g2846 (n2040, n479, n_1204);
  not g2851 (n_1207, n2042);
  and g2852 (n2043, n_182, n_1207);
  and g2853 (n2044, n275, n_305);
  and g2854 (n2045, n288, n_296);
  and g2858 (n2047, n302, n_326);
  and g2859 (n2048, n315, n_317);
  not g2864 (n_1212, n2050);
  and g2865 (n2051, n479, n_1212);
  and g2866 (n2052, n275, n_46);
  and g2867 (n2053, n288, n_37);
  and g2871 (n2055, n302, n_285);
  and g2872 (n2056, n315, n_276);
  not g2877 (n_1217, n2058);
  and g2878 (n2059, n426, n_1217);
  and g2882 (n2061, n275, n_346);
  and g2883 (n2062, n288, n_337);
  and g2887 (n2064, n302, n_242);
  and g2888 (n2065, n315, n_233);
  not g2893 (n_1224, n2067);
  and g2894 (n2068, n372, n_1224);
  and g2895 (n2069, n275, n_262);
  and g2896 (n2070, n288, n_253);
  and g2900 (n2072, n302, n_201);
  and g2901 (n2073, n315, n_192);
  not g2906 (n_1229, n2075);
  and g2907 (n2076, n319, n_1229);
  not g2912 (n_1232, n2078);
  and g2913 (n2079, \shift[6] , n_1232);
  or g2914 (\result[8] , n2043, n2079);
  and g2915 (n2081, n275, n_399);
  and g2916 (n2082, n288, n_394);
  and g2920 (n2084, n302, n_362);
  and g2921 (n2085, n315, n_357);
  not g2926 (n_1237, n2087);
  and g2927 (n2088, n319, n_1237);
  and g2928 (n2089, n275, n_451);
  and g2929 (n2090, n288, n_446);
  and g2933 (n2092, n302, n_387);
  and g2934 (n2093, n315, n_382);
  not g2939 (n_1242, n2095);
  and g2940 (n2096, n372, n_1242);
  and g2944 (n2098, n275, n_504);
  and g2945 (n2099, n288, n_499);
  and g2949 (n2101, n302, n_414);
  and g2950 (n2102, n315, n_409);
  not g2955 (n_1249, n2104);
  and g2956 (n2105, n426, n_1249);
  and g2957 (n2106, n275, n_426);
  and g2958 (n2107, n288, n_421);
  and g2962 (n2109, n302, n_439);
  and g2963 (n2110, n315, n_434);
  not g2968 (n_1254, n2112);
  and g2969 (n2113, n479, n_1254);
  not g2974 (n_1257, n2115);
  and g2975 (n2116, n_182, n_1257);
  and g2976 (n2117, n275, n_479);
  and g2977 (n2118, n288, n_474);
  and g2981 (n2120, n302, n_519);
  and g2982 (n2121, n315, n_514);
  not g2987 (n_1262, n2123);
  and g2988 (n2124, n479, n_1262);
  and g2989 (n2125, n275, n_374);
  and g2990 (n2126, n288, n_369);
  and g2994 (n2128, n302, n_467);
  and g2995 (n2129, n315, n_462);
  not g3000 (n_1267, n2131);
  and g3001 (n2132, n426, n_1267);
  and g3005 (n2134, n275, n_531);
  and g3006 (n2135, n288, n_526);
  and g3010 (n2137, n302, n_544);
  and g3011 (n2138, n315, n_539);
  not g3016 (n_1274, n2140);
  and g3017 (n2141, n372, n_1274);
  and g3018 (n2142, n275, n_556);
  and g3019 (n2143, n288, n_551);
  and g3023 (n2145, n302, n_492);
  and g3024 (n2146, n315, n_487);
  not g3029 (n_1279, n2148);
  and g3030 (n2149, n319, n_1279);
  not g3035 (n_1282, n2151);
  and g3036 (n2152, \shift[6] , n_1282);
  or g3037 (\result[9] , n2116, n2152);
  and g3038 (n2154, n275, n_609);
  and g3039 (n2155, n288, n_604);
  and g3043 (n2157, n302, n_572);
  and g3044 (n2158, n315, n_567);
  not g3049 (n_1287, n2160);
  and g3050 (n2161, n319, n_1287);
  and g3051 (n2162, n275, n_661);
  and g3052 (n2163, n288, n_656);
  and g3056 (n2165, n302, n_597);
  and g3057 (n2166, n315, n_592);
  not g3062 (n_1292, n2168);
  and g3063 (n2169, n372, n_1292);
  and g3067 (n2171, n275, n_714);
  and g3068 (n2172, n288, n_709);
  and g3072 (n2174, n302, n_624);
  and g3073 (n2175, n315, n_619);
  not g3078 (n_1299, n2177);
  and g3079 (n2178, n426, n_1299);
  and g3080 (n2179, n275, n_636);
  and g3081 (n2180, n288, n_631);
  and g3085 (n2182, n302, n_649);
  and g3086 (n2183, n315, n_644);
  not g3091 (n_1304, n2185);
  and g3092 (n2186, n479, n_1304);
  not g3097 (n_1307, n2188);
  and g3098 (n2189, n_182, n_1307);
  and g3099 (n2190, n275, n_689);
  and g3100 (n2191, n288, n_684);
  and g3104 (n2193, n302, n_729);
  and g3105 (n2194, n315, n_724);
  not g3110 (n_1312, n2196);
  and g3111 (n2197, n479, n_1312);
  and g3112 (n2198, n275, n_584);
  and g3113 (n2199, n288, n_579);
  and g3117 (n2201, n302, n_677);
  and g3118 (n2202, n315, n_672);
  not g3123 (n_1317, n2204);
  and g3124 (n2205, n426, n_1317);
  and g3128 (n2207, n275, n_741);
  and g3129 (n2208, n288, n_736);
  and g3133 (n2210, n302, n_754);
  and g3134 (n2211, n315, n_749);
  not g3139 (n_1324, n2213);
  and g3140 (n2214, n372, n_1324);
  and g3141 (n2215, n275, n_766);
  and g3142 (n2216, n288, n_761);
  and g3146 (n2218, n302, n_702);
  and g3147 (n2219, n315, n_697);
  not g3152 (n_1329, n2221);
  and g3153 (n2222, n319, n_1329);
  not g3158 (n_1332, n2224);
  and g3159 (n2225, \shift[6] , n_1332);
  or g3160 (\result[10] , n2189, n2225);
  and g3161 (n2227, n275, n_819);
  and g3162 (n2228, n288, n_814);
  and g3166 (n2230, n302, n_859);
  and g3167 (n2231, n315, n_854);
  not g3172 (n_1337, n2233);
  and g3173 (n2234, n319, n_1337);
  and g3174 (n2235, n275, n_794);
  and g3175 (n2236, n288, n_789);
  and g3179 (n2238, n302, n_807);
  and g3180 (n2239, n315, n_802);
  not g3185 (n_1342, n2241);
  and g3186 (n2242, n372, n_1342);
  and g3190 (n2244, n275, n_951);
  and g3191 (n2245, n288, n_946);
  and g3195 (n2247, n302, n_834);
  and g3196 (n2248, n315, n_829);
  not g3201 (n_1349, n2250);
  and g3202 (n2251, n426, n_1349);
  and g3203 (n2252, n275, n_846);
  and g3204 (n2253, n288, n_841);
  and g3208 (n2255, n302, n_782);
  and g3209 (n2256, n315, n_777);
  not g3214 (n_1354, n2258);
  and g3215 (n2259, n479, n_1354);
  not g3220 (n_1357, n2261);
  and g3221 (n2262, n_182, n_1357);
  and g3222 (n2263, n275, n_899);
  and g3223 (n2264, n315, n_907);
  and g3227 (n2266, n302, n_912);
  and g3228 (n2267, n288, n_894);
  not g3233 (n_1362, n2269);
  and g3234 (n2270, n479, n_1362);
  and g3235 (n2271, n275, n_871);
  and g3236 (n2272, n288, n_866);
  and g3240 (n2274, n302, n_887);
  and g3241 (n2275, n315, n_882);
  not g3246 (n_1367, n2277);
  and g3247 (n2278, n426, n_1367);
  and g3251 (n2280, n275, n_924);
  and g3252 (n2281, n288, n_919);
  and g3256 (n2283, n302, n_964);
  and g3257 (n2284, n315, n_959);
  not g3262 (n_1374, n2286);
  and g3263 (n2287, n372, n_1374);
  and g3264 (n2288, n275, n_976);
  and g3265 (n2289, n288, n_971);
  and g3269 (n2291, n302, n_939);
  and g3270 (n2292, n315, n_934);
  not g3275 (n_1379, n2294);
  and g3276 (n2295, n319, n_1379);
  not g3281 (n_1382, n2297);
  and g3282 (n2298, \shift[6] , n_1382);
  or g3283 (\result[11] , n2262, n2298);
  and g3284 (n2300, n275, n_69);
  and g3285 (n2301, n288, n_89);
  and g3289 (n2303, n_17, n302);
  and g3290 (n2304, n315, n_80);
  not g3295 (n_1387, n2306);
  and g3296 (n2307, n319, n_1387);
  and g3297 (n2308, n275, n_155);
  and g3298 (n2309, n288, n_175);
  and g3302 (n2311, n302, n_60);
  and g3303 (n2312, n315, n_166);
  not g3308 (n_1392, n2314);
  and g3309 (n2315, n372, n_1392);
  and g3313 (n2317, n275, n_201);
  and g3314 (n2318, n288, n_221);
  and g3318 (n2320, n302, n_104);
  and g3319 (n2321, n315, n_212);
  not g3324 (n_1399, n2323);
  and g3325 (n2324, n426, n_1399);
  and g3326 (n2325, n275, n_113);
  and g3327 (n2326, n288, n_133);
  and g3331 (n2328, n302, n_146);
  and g3332 (n2329, n315, n_124);
  not g3337 (n_1404, n2331);
  and g3338 (n2332, n479, n_1404);
  not g3343 (n_1407, n2334);
  and g3344 (n2335, n_182, n_1407);
  and g3345 (n2336, n275, n_285);
  and g3346 (n2337, n288, n_305);
  and g3350 (n2339, n302, n_317);
  and g3351 (n2340, n315, n_296);
  not g3356 (n_1412, n2342);
  and g3357 (n2343, n479, n_1412);
  and g3358 (n2344, n275, n_26);
  and g3359 (n2345, n288, n_46);
  and g3363 (n2347, n302, n_276);
  and g3364 (n2348, n_37, n315);
  not g3369 (n_1417, n2350);
  and g3370 (n2351, n426, n_1417);
  and g3374 (n2353, n275, n_326);
  and g3375 (n2354, n288, n_346);
  and g3379 (n2356, n302, n_233);
  and g3380 (n2357, n315, n_337);
  not g3385 (n_1424, n2359);
  and g3386 (n2360, n372, n_1424);
  and g3387 (n2361, n275, n_242);
  and g3388 (n2362, n288, n_262);
  and g3392 (n2364, n302, n_192);
  and g3393 (n2365, n315, n_253);
  not g3398 (n_1429, n2367);
  and g3399 (n2368, n319, n_1429);
  not g3404 (n_1432, n2370);
  and g3405 (n2371, \shift[6] , n_1432);
  or g3406 (\result[12] , n2335, n2371);
  and g3407 (n2373, n275, n_387);
  and g3408 (n2374, n288, n_399);
  and g3412 (n2376, n302, n_357);
  and g3413 (n2377, n315, n_394);
  not g3418 (n_1437, n2379);
  and g3419 (n2380, n319, n_1437);
  and g3420 (n2381, n275, n_439);
  and g3421 (n2382, n288, n_451);
  and g3425 (n2384, n302, n_382);
  and g3426 (n2385, n315, n_446);
  not g3431 (n_1442, n2387);
  and g3432 (n2388, n372, n_1442);
  and g3436 (n2390, n275, n_492);
  and g3437 (n2391, n288, n_504);
  and g3441 (n2393, n302, n_409);
  and g3442 (n2394, n315, n_499);
  not g3447 (n_1449, n2396);
  and g3448 (n2397, n426, n_1449);
  and g3449 (n2398, n275, n_414);
  and g3450 (n2399, n288, n_426);
  and g3454 (n2401, n302, n_434);
  and g3455 (n2402, n315, n_421);
  not g3460 (n_1454, n2404);
  and g3461 (n2405, n479, n_1454);
  not g3466 (n_1457, n2407);
  and g3467 (n2408, n_182, n_1457);
  and g3468 (n2409, n275, n_467);
  and g3469 (n2410, n288, n_479);
  and g3473 (n2412, n302, n_514);
  and g3474 (n2413, n315, n_474);
  not g3479 (n_1462, n2415);
  and g3480 (n2416, n479, n_1462);
  and g3481 (n2417, n275, n_362);
  and g3482 (n2418, n288, n_374);
  and g3486 (n2420, n302, n_462);
  and g3487 (n2421, n315, n_369);
  not g3492 (n_1467, n2423);
  and g3493 (n2424, n426, n_1467);
  and g3497 (n2426, n275, n_519);
  and g3498 (n2427, n288, n_531);
  and g3502 (n2429, n302, n_539);
  and g3503 (n2430, n315, n_526);
  not g3508 (n_1474, n2432);
  and g3509 (n2433, n372, n_1474);
  and g3510 (n2434, n275, n_544);
  and g3511 (n2435, n288, n_556);
  and g3515 (n2437, n302, n_487);
  and g3516 (n2438, n315, n_551);
  not g3521 (n_1479, n2440);
  and g3522 (n2441, n319, n_1479);
  not g3527 (n_1482, n2443);
  and g3528 (n2444, \shift[6] , n_1482);
  or g3529 (\result[13] , n2408, n2444);
  and g3530 (n2446, n275, n_597);
  and g3531 (n2447, n288, n_609);
  and g3535 (n2449, n302, n_567);
  and g3536 (n2450, n315, n_604);
  not g3541 (n_1487, n2452);
  and g3542 (n2453, n319, n_1487);
  and g3543 (n2454, n275, n_649);
  and g3544 (n2455, n288, n_661);
  and g3548 (n2457, n302, n_592);
  and g3549 (n2458, n315, n_656);
  not g3554 (n_1492, n2460);
  and g3555 (n2461, n372, n_1492);
  and g3559 (n2463, n275, n_702);
  and g3560 (n2464, n288, n_714);
  and g3564 (n2466, n302, n_619);
  and g3565 (n2467, n315, n_709);
  not g3570 (n_1499, n2469);
  and g3571 (n2470, n426, n_1499);
  and g3572 (n2471, n275, n_624);
  and g3573 (n2472, n288, n_636);
  and g3577 (n2474, n302, n_644);
  and g3578 (n2475, n315, n_631);
  not g3583 (n_1504, n2477);
  and g3584 (n2478, n479, n_1504);
  not g3589 (n_1507, n2480);
  and g3590 (n2481, n_182, n_1507);
  and g3591 (n2482, n275, n_677);
  and g3592 (n2483, n288, n_689);
  and g3596 (n2485, n302, n_724);
  and g3597 (n2486, n315, n_684);
  not g3602 (n_1512, n2488);
  and g3603 (n2489, n479, n_1512);
  and g3604 (n2490, n275, n_572);
  and g3605 (n2491, n288, n_584);
  and g3609 (n2493, n302, n_672);
  and g3610 (n2494, n315, n_579);
  not g3615 (n_1517, n2496);
  and g3616 (n2497, n426, n_1517);
  and g3620 (n2499, n275, n_729);
  and g3621 (n2500, n288, n_741);
  and g3625 (n2502, n302, n_749);
  and g3626 (n2503, n315, n_736);
  not g3631 (n_1524, n2505);
  and g3632 (n2506, n372, n_1524);
  and g3633 (n2507, n275, n_754);
  and g3634 (n2508, n288, n_766);
  and g3638 (n2510, n302, n_697);
  and g3639 (n2511, n315, n_761);
  not g3644 (n_1529, n2513);
  and g3645 (n2514, n319, n_1529);
  not g3650 (n_1532, n2516);
  and g3651 (n2517, \shift[6] , n_1532);
  or g3652 (\result[14] , n2481, n2517);
  and g3653 (n2519, n275, n_807);
  and g3654 (n2520, n288, n_819);
  and g3658 (n2522, n302, n_854);
  and g3659 (n2523, n315, n_814);
  not g3664 (n_1537, n2525);
  and g3665 (n2526, n319, n_1537);
  and g3666 (n2527, n275, n_782);
  and g3667 (n2528, n288, n_794);
  and g3671 (n2530, n302, n_802);
  and g3672 (n2531, n315, n_789);
  not g3677 (n_1542, n2533);
  and g3678 (n2534, n372, n_1542);
  and g3682 (n2536, n275, n_939);
  and g3683 (n2537, n288, n_951);
  and g3687 (n2539, n302, n_829);
  and g3688 (n2540, n315, n_946);
  not g3693 (n_1549, n2542);
  and g3694 (n2543, n426, n_1549);
  and g3695 (n2544, n275, n_834);
  and g3696 (n2545, n288, n_846);
  and g3700 (n2547, n302, n_777);
  and g3701 (n2548, n315, n_841);
  not g3706 (n_1554, n2550);
  and g3707 (n2551, n479, n_1554);
  not g3712 (n_1557, n2553);
  and g3713 (n2554, n_182, n_1557);
  and g3714 (n2555, n275, n_887);
  and g3715 (n2556, n288, n_899);
  and g3719 (n2558, n302, n_907);
  and g3720 (n2559, n315, n_894);
  not g3725 (n_1562, n2561);
  and g3726 (n2562, n479, n_1562);
  and g3727 (n2563, n275, n_859);
  and g3728 (n2564, n288, n_871);
  and g3732 (n2566, n302, n_882);
  and g3733 (n2567, n315, n_866);
  not g3738 (n_1567, n2569);
  and g3739 (n2570, n426, n_1567);
  and g3743 (n2572, n275, n_912);
  and g3744 (n2573, n288, n_924);
  and g3748 (n2575, n302, n_959);
  and g3749 (n2576, n315, n_919);
  not g3754 (n_1574, n2578);
  and g3755 (n2579, n372, n_1574);
  and g3756 (n2580, n275, n_964);
  and g3757 (n2581, n288, n_976);
  and g3761 (n2583, n302, n_934);
  and g3762 (n2584, n315, n_971);
  not g3767 (n_1579, n2586);
  and g3768 (n2587, n319, n_1579);
  not g3773 (n_1582, n2589);
  and g3774 (n2590, \shift[6] , n_1582);
  or g3775 (\result[15] , n2554, n2590);
  and g3776 (n2592, n319, n_93);
  and g3777 (n2593, n372, n_178);
  and g3781 (n2595, n426, n_224);
  and g3782 (n2596, n_137, n479);
  not g3787 (n_1587, n2598);
  and g3788 (n2599, n_182, n_1587);
  and g3789 (n2600, n_51, n426);
  and g3790 (n2601, n319, n_265);
  and g3794 (n2603, n479, n_308);
  and g3795 (n2604, n372, n_349);
  not g3800 (n_1592, n2606);
  and g3801 (n2607, \shift[6] , n_1592);
  or g3802 (\result[16] , n2599, n2607);
  and g3803 (n2609, n319, n_402);
  and g3804 (n2610, n372, n_454);
  and g3808 (n2612, n426, n_507);
  and g3809 (n2613, n479, n_429);
  not g3814 (n_1597, n2615);
  and g3815 (n2616, n_182, n_1597);
  and g3816 (n2617, n479, n_482);
  and g3817 (n2618, n426, n_377);
  and g3821 (n2620, n372, n_534);
  and g3822 (n2621, n319, n_559);
  not g3827 (n_1602, n2623);
  and g3828 (n2624, \shift[6] , n_1602);
  or g3829 (\result[17] , n2616, n2624);
  and g3830 (n2626, n319, n_612);
  and g3831 (n2627, n372, n_664);
  and g3835 (n2629, n426, n_717);
  and g3836 (n2630, n479, n_639);
  not g3841 (n_1607, n2632);
  and g3842 (n2633, n_182, n_1607);
  and g3843 (n2634, n479, n_692);
  and g3844 (n2635, n426, n_587);
  and g3848 (n2637, n372, n_744);
  and g3849 (n2638, n319, n_769);
  not g3854 (n_1612, n2640);
  and g3855 (n2641, \shift[6] , n_1612);
  or g3856 (\result[18] , n2633, n2641);
  and g3857 (n2643, n372, n_797);
  and g3858 (n2644, n319, n_822);
  and g3862 (n2646, n479, n_849);
  and g3863 (n2647, n426, n_954);
  not g3868 (n_1617, n2649);
  and g3869 (n2650, n_182, n_1617);
  and g3870 (n2651, n479, n_902);
  and g3871 (n2652, n426, n_874);
  and g3875 (n2654, n319, n_979);
  and g3876 (n2655, n372, n_927);
  not g3881 (n_1622, n2657);
  and g3882 (n2658, \shift[6] , n_1622);
  or g3883 (\result[19] , n2650, n2658);
  and g3884 (n2660, n319, n_992);
  and g3885 (n2661, n372, n_1004);
  and g3889 (n2663, n426, n_1029);
  and g3890 (n2664, n479, n_999);
  not g3895 (n_1627, n2666);
  and g3896 (n2667, n_182, n_1627);
  and g3897 (n2668, n426, n_987);
  and g3898 (n2669, n372, n_1012);
  and g3902 (n2671, n319, n_1024);
  and g3903 (n2672, n479, n_1017);
  not g3908 (n_1632, n2674);
  and g3909 (n2675, \shift[6] , n_1632);
  or g3910 (\result[20] , n2667, n2675);
  and g3911 (n2677, n319, n_1042);
  and g3912 (n2678, n372, n_1054);
  and g3916 (n2680, n426, n_1079);
  and g3917 (n2681, n479, n_1049);
  not g3922 (n_1637, n2683);
  and g3923 (n2684, n_182, n_1637);
  and g3924 (n2685, n426, n_1037);
  and g3925 (n2686, n372, n_1062);
  and g3929 (n2688, n319, n_1074);
  and g3930 (n2689, n479, n_1067);
  not g3935 (n_1642, n2691);
  and g3936 (n2692, \shift[6] , n_1642);
  or g3937 (\result[21] , n2684, n2692);
  and g3938 (n2694, n319, n_1092);
  and g3939 (n2695, n372, n_1104);
  and g3943 (n2697, n426, n_1129);
  and g3944 (n2698, n479, n_1099);
  not g3949 (n_1647, n2700);
  and g3950 (n2701, n_182, n_1647);
  and g3951 (n2702, n426, n_1087);
  and g3952 (n2703, n372, n_1112);
  and g3956 (n2705, n319, n_1124);
  and g3957 (n2706, n479, n_1117);
  not g3962 (n_1652, n2708);
  and g3963 (n2709, \shift[6] , n_1652);
  or g3964 (\result[22] , n2701, n2709);
  and g3965 (n2711, n319, n_1142);
  and g3966 (n2712, n426, n_1179);
  and g3970 (n2714, n479, n_1149);
  and g3971 (n2715, n372, n_1154);
  not g3976 (n_1657, n2717);
  and g3977 (n2718, n_182, n_1657);
  and g3978 (n2719, n372, n_1162);
  and g3979 (n2720, n479, n_1167);
  and g3983 (n2722, n319, n_1174);
  and g3984 (n2723, n426, n_1137);
  not g3989 (n_1662, n2725);
  and g3990 (n2726, \shift[6] , n_1662);
  or g3991 (\result[23] , n2718, n2726);
  and g3992 (n2728, n319, n_1192);
  and g3993 (n2729, n426, n_1229);
  and g3997 (n2731, n479, n_1199);
  and g3998 (n2732, n372, n_1204);
  not g4003 (n_1667, n2734);
  and g4004 (n2735, n_182, n_1667);
  and g4005 (n2736, n372, n_1212);
  and g4006 (n2737, n479, n_1217);
  and g4010 (n2739, n319, n_1224);
  and g4011 (n2740, n426, n_1187);
  not g4016 (n_1672, n2742);
  and g4017 (n2743, \shift[6] , n_1672);
  or g4018 (\result[24] , n2735, n2743);
  and g4019 (n2745, n319, n_1242);
  and g4020 (n2746, n426, n_1279);
  and g4024 (n2748, n479, n_1249);
  and g4025 (n2749, n372, n_1254);
  not g4030 (n_1677, n2751);
  and g4031 (n2752, n_182, n_1677);
  and g4032 (n2753, n372, n_1262);
  and g4033 (n2754, n479, n_1267);
  and g4037 (n2756, n319, n_1274);
  and g4038 (n2757, n426, n_1237);
  not g4043 (n_1682, n2759);
  and g4044 (n2760, \shift[6] , n_1682);
  or g4045 (\result[25] , n2752, n2760);
  and g4046 (n2762, n319, n_1292);
  and g4047 (n2763, n372, n_1304);
  and g4051 (n2765, n426, n_1329);
  and g4052 (n2766, n479, n_1299);
  not g4057 (n_1687, n2768);
  and g4058 (n2769, n_182, n_1687);
  and g4059 (n2770, n372, n_1312);
  and g4060 (n2771, n479, n_1317);
  and g4064 (n2773, n319, n_1324);
  and g4065 (n2774, n426, n_1287);
  not g4070 (n_1692, n2776);
  and g4071 (n2777, \shift[6] , n_1692);
  or g4072 (\result[26] , n2769, n2777);
  and g4073 (n2779, n319, n_1342);
  and g4074 (n2780, n372, n_1354);
  and g4078 (n2782, n426, n_1379);
  and g4079 (n2783, n479, n_1349);
  not g4084 (n_1697, n2785);
  and g4085 (n2786, n_182, n_1697);
  and g4086 (n2787, n372, n_1362);
  and g4087 (n2788, n479, n_1367);
  and g4091 (n2790, n319, n_1374);
  and g4092 (n2791, n426, n_1337);
  not g4097 (n_1702, n2793);
  and g4098 (n2794, \shift[6] , n_1702);
  or g4099 (\result[27] , n2786, n2794);
  and g4100 (n2796, n319, n_1392);
  and g4101 (n2797, n372, n_1404);
  and g4105 (n2799, n426, n_1429);
  and g4106 (n2800, n479, n_1399);
  not g4111 (n_1707, n2802);
  and g4112 (n2803, n_182, n_1707);
  and g4113 (n2804, n372, n_1412);
  and g4114 (n2805, n479, n_1417);
  and g4118 (n2807, n319, n_1424);
  and g4119 (n2808, n426, n_1387);
  not g4124 (n_1712, n2810);
  and g4125 (n2811, \shift[6] , n_1712);
  or g4126 (\result[28] , n2803, n2811);
  and g4127 (n2813, n319, n_1442);
  and g4128 (n2814, n372, n_1454);
  and g4132 (n2816, n426, n_1479);
  and g4133 (n2817, n479, n_1449);
  not g4138 (n_1717, n2819);
  and g4139 (n2820, n_182, n_1717);
  and g4140 (n2821, n372, n_1462);
  and g4141 (n2822, n479, n_1467);
  and g4145 (n2824, n319, n_1474);
  and g4146 (n2825, n426, n_1437);
  not g4151 (n_1722, n2827);
  and g4152 (n2828, \shift[6] , n_1722);
  or g4153 (\result[29] , n2820, n2828);
  and g4154 (n2830, n319, n_1492);
  and g4155 (n2831, n372, n_1504);
  and g4159 (n2833, n426, n_1529);
  and g4160 (n2834, n479, n_1499);
  not g4165 (n_1727, n2836);
  and g4166 (n2837, n_182, n_1727);
  and g4167 (n2838, n372, n_1512);
  and g4168 (n2839, n479, n_1517);
  and g4172 (n2841, n319, n_1524);
  and g4173 (n2842, n426, n_1487);
  not g4178 (n_1732, n2844);
  and g4179 (n2845, \shift[6] , n_1732);
  or g4180 (\result[30] , n2837, n2845);
  and g4181 (n2847, n319, n_1542);
  and g4182 (n2848, n372, n_1554);
  and g4186 (n2850, n426, n_1579);
  and g4187 (n2851, n479, n_1549);
  not g4192 (n_1737, n2853);
  and g4193 (n2854, n_182, n_1737);
  and g4194 (n2855, n372, n_1562);
  and g4195 (n2856, n479, n_1567);
  and g4199 (n2858, n319, n_1574);
  and g4200 (n2859, n426, n_1537);
  not g4205 (n_1742, n2861);
  and g4206 (n2862, \shift[6] , n_1742);
  or g4207 (\result[31] , n2854, n2862);
  and g4208 (n2864, n319, n_178);
  and g4209 (n2865, n372, n_137);
  and g4213 (n2867, n426, n_265);
  and g4214 (n2868, n479, n_224);
  not g4219 (n_1747, n2870);
  and g4220 (n2871, n_182, n_1747);
  and g4221 (n2872, n_51, n479);
  and g4222 (n2873, n_93, n426);
  and g4226 (n2875, n372, n_308);
  and g4227 (n2876, n319, n_349);
  not g4232 (n_1752, n2878);
  and g4233 (n2879, \shift[6] , n_1752);
  or g4234 (\result[32] , n2871, n2879);
  and g4235 (n2881, n319, n_454);
  and g4236 (n2882, n372, n_429);
  and g4240 (n2884, n426, n_559);
  and g4241 (n2885, n479, n_507);
  not g4246 (n_1757, n2887);
  and g4247 (n2888, n_182, n_1757);
  and g4248 (n2889, n372, n_482);
  and g4249 (n2890, n479, n_377);
  and g4253 (n2892, n319, n_534);
  and g4254 (n2893, n426, n_402);
  not g4259 (n_1762, n2895);
  and g4260 (n2896, \shift[6] , n_1762);
  or g4261 (\result[33] , n2888, n2896);
  and g4262 (n2898, n319, n_664);
  and g4263 (n2899, n372, n_639);
  and g4267 (n2901, n426, n_769);
  and g4268 (n2902, n479, n_717);
  not g4273 (n_1767, n2904);
  and g4274 (n2905, n_182, n_1767);
  and g4275 (n2906, n372, n_692);
  and g4276 (n2907, n479, n_587);
  and g4280 (n2909, n319, n_744);
  and g4281 (n2910, n426, n_612);
  not g4286 (n_1772, n2912);
  and g4287 (n2913, \shift[6] , n_1772);
  or g4288 (\result[34] , n2905, n2913);
  and g4289 (n2915, n319, n_797);
  and g4290 (n2916, n426, n_979);
  and g4294 (n2918, n372, n_849);
  and g4295 (n2919, n479, n_954);
  not g4300 (n_1777, n2921);
  and g4301 (n2922, n_182, n_1777);
  and g4302 (n2923, n372, n_902);
  and g4303 (n2924, n426, n_822);
  and g4307 (n2926, n319, n_927);
  and g4308 (n2927, n479, n_874);
  not g4313 (n_1782, n2929);
  and g4314 (n2930, \shift[6] , n_1782);
  or g4315 (\result[35] , n2922, n2930);
  and g4316 (n2932, n319, n_1004);
  and g4317 (n2933, n372, n_999);
  and g4321 (n2935, n426, n_1024);
  and g4322 (n2936, n479, n_1029);
  not g4327 (n_1787, n2938);
  and g4328 (n2939, n_182, n_1787);
  and g4329 (n2940, n479, n_987);
  and g4330 (n2941, n426, n_992);
  and g4334 (n2943, n372, n_1017);
  and g4335 (n2944, n319, n_1012);
  not g4340 (n_1792, n2946);
  and g4341 (n2947, \shift[6] , n_1792);
  or g4342 (\result[36] , n2939, n2947);
  and g4343 (n2949, n319, n_1054);
  and g4344 (n2950, n372, n_1049);
  and g4348 (n2952, n426, n_1074);
  and g4349 (n2953, n479, n_1079);
  not g4354 (n_1797, n2955);
  and g4355 (n2956, n_182, n_1797);
  and g4356 (n2957, n479, n_1037);
  and g4357 (n2958, n426, n_1042);
  and g4361 (n2960, n372, n_1067);
  and g4362 (n2961, n319, n_1062);
  not g4367 (n_1802, n2963);
  and g4368 (n2964, \shift[6] , n_1802);
  or g4369 (\result[37] , n2956, n2964);
  and g4370 (n2966, n319, n_1104);
  and g4371 (n2967, n372, n_1099);
  and g4375 (n2969, n426, n_1124);
  and g4376 (n2970, n479, n_1129);
  not g4381 (n_1807, n2972);
  and g4382 (n2973, n_182, n_1807);
  and g4383 (n2974, n479, n_1087);
  and g4384 (n2975, n426, n_1092);
  and g4388 (n2977, n372, n_1117);
  and g4389 (n2978, n319, n_1112);
  not g4394 (n_1812, n2980);
  and g4395 (n2981, \shift[6] , n_1812);
  or g4396 (\result[38] , n2973, n2981);
  and g4397 (n2983, n479, n_1179);
  and g4398 (n2984, n426, n_1174);
  and g4402 (n2986, n372, n_1149);
  and g4403 (n2987, n319, n_1154);
  not g4408 (n_1817, n2989);
  and g4409 (n2990, n_182, n_1817);
  and g4410 (n2991, n319, n_1162);
  and g4411 (n2992, n372, n_1167);
  and g4415 (n2994, n426, n_1142);
  and g4416 (n2995, n479, n_1137);
  not g4421 (n_1822, n2997);
  and g4422 (n2998, \shift[6] , n_1822);
  or g4423 (\result[39] , n2990, n2998);
  and g4424 (n3000, n479, n_1229);
  and g4425 (n3001, n426, n_1224);
  and g4429 (n3003, n372, n_1199);
  and g4430 (n3004, n319, n_1204);
  not g4435 (n_1827, n3006);
  and g4436 (n3007, n_182, n_1827);
  and g4437 (n3008, n319, n_1212);
  and g4438 (n3009, n372, n_1217);
  and g4442 (n3011, n426, n_1192);
  and g4443 (n3012, n479, n_1187);
  not g4448 (n_1832, n3014);
  and g4449 (n3015, \shift[6] , n_1832);
  or g4450 (\result[40] , n3007, n3015);
  and g4451 (n3017, n479, n_1279);
  and g4452 (n3018, n426, n_1274);
  and g4456 (n3020, n372, n_1249);
  and g4457 (n3021, n319, n_1254);
  not g4462 (n_1837, n3023);
  and g4463 (n3024, n_182, n_1837);
  and g4464 (n3025, n319, n_1262);
  and g4465 (n3026, n372, n_1267);
  and g4469 (n3028, n426, n_1242);
  and g4470 (n3029, n479, n_1237);
  not g4475 (n_1842, n3031);
  and g4476 (n3032, \shift[6] , n_1842);
  or g4477 (\result[41] , n3024, n3032);
  and g4478 (n3034, n319, n_1304);
  and g4479 (n3035, n372, n_1299);
  and g4483 (n3037, n426, n_1324);
  and g4484 (n3038, n479, n_1329);
  not g4489 (n_1847, n3040);
  and g4490 (n3041, n_182, n_1847);
  and g4491 (n3042, n319, n_1312);
  and g4492 (n3043, n372, n_1317);
  and g4496 (n3045, n426, n_1292);
  and g4497 (n3046, n479, n_1287);
  not g4502 (n_1852, n3048);
  and g4503 (n3049, \shift[6] , n_1852);
  or g4504 (\result[42] , n3041, n3049);
  and g4505 (n3051, n319, n_1354);
  and g4506 (n3052, n372, n_1349);
  and g4510 (n3054, n426, n_1374);
  and g4511 (n3055, n479, n_1379);
  not g4516 (n_1857, n3057);
  and g4517 (n3058, n_182, n_1857);
  and g4518 (n3059, n319, n_1362);
  and g4519 (n3060, n372, n_1367);
  and g4523 (n3062, n426, n_1342);
  and g4524 (n3063, n479, n_1337);
  not g4529 (n_1862, n3065);
  and g4530 (n3066, \shift[6] , n_1862);
  or g4531 (\result[43] , n3058, n3066);
  and g4532 (n3068, n319, n_1404);
  and g4533 (n3069, n372, n_1399);
  and g4537 (n3071, n426, n_1424);
  and g4538 (n3072, n479, n_1429);
  not g4543 (n_1867, n3074);
  and g4544 (n3075, n_182, n_1867);
  and g4545 (n3076, n319, n_1412);
  and g4546 (n3077, n372, n_1417);
  and g4550 (n3079, n426, n_1392);
  and g4551 (n3080, n479, n_1387);
  not g4556 (n_1872, n3082);
  and g4557 (n3083, \shift[6] , n_1872);
  or g4558 (\result[44] , n3075, n3083);
  and g4559 (n3085, n319, n_1454);
  and g4560 (n3086, n372, n_1449);
  and g4564 (n3088, n426, n_1474);
  and g4565 (n3089, n479, n_1479);
  not g4570 (n_1877, n3091);
  and g4571 (n3092, n_182, n_1877);
  and g4572 (n3093, n319, n_1462);
  and g4573 (n3094, n372, n_1467);
  and g4577 (n3096, n426, n_1442);
  and g4578 (n3097, n479, n_1437);
  not g4583 (n_1882, n3099);
  and g4584 (n3100, \shift[6] , n_1882);
  or g4585 (\result[45] , n3092, n3100);
  and g4586 (n3102, n319, n_1504);
  and g4587 (n3103, n372, n_1499);
  and g4591 (n3105, n426, n_1524);
  and g4592 (n3106, n479, n_1529);
  not g4597 (n_1887, n3108);
  and g4598 (n3109, n_182, n_1887);
  and g4599 (n3110, n319, n_1512);
  and g4600 (n3111, n372, n_1517);
  and g4604 (n3113, n426, n_1492);
  and g4605 (n3114, n479, n_1487);
  not g4610 (n_1892, n3116);
  and g4611 (n3117, \shift[6] , n_1892);
  or g4612 (\result[46] , n3109, n3117);
  and g4613 (n3119, n319, n_1554);
  and g4614 (n3120, n372, n_1549);
  and g4618 (n3122, n426, n_1574);
  and g4619 (n3123, n479, n_1579);
  not g4624 (n_1897, n3125);
  and g4625 (n3126, n_182, n_1897);
  and g4626 (n3127, n319, n_1562);
  and g4627 (n3128, n372, n_1567);
  and g4631 (n3130, n426, n_1542);
  and g4632 (n3131, n479, n_1537);
  not g4637 (n_1902, n3133);
  and g4638 (n3134, \shift[6] , n_1902);
  or g4639 (\result[47] , n3126, n3134);
  and g4640 (n3136, n319, n_137);
  and g4641 (n3137, n372, n_224);
  and g4645 (n3139, n426, n_349);
  and g4646 (n3140, n479, n_265);
  not g4651 (n_1907, n3142);
  and g4652 (n3143, n_182, n_1907);
  and g4653 (n3144, n_51, n372);
  and g4654 (n3145, n_93, n479);
  and g4658 (n3147, n319, n_308);
  and g4659 (n3148, n426, n_178);
  not g4664 (n_1912, n3150);
  and g4665 (n3151, \shift[6] , n_1912);
  or g4666 (\result[48] , n3143, n3151);
  and g4667 (n3153, n319, n_429);
  and g4668 (n3154, n372, n_507);
  and g4672 (n3156, n426, n_534);
  and g4673 (n3157, n479, n_559);
  not g4678 (n_1917, n3159);
  and g4679 (n3160, n_182, n_1917);
  and g4680 (n3161, n319, n_482);
  and g4681 (n3162, n372, n_377);
  and g4685 (n3164, n426, n_454);
  and g4686 (n3165, n479, n_402);
  not g4691 (n_1922, n3167);
  and g4692 (n3168, \shift[6] , n_1922);
  or g4693 (\result[49] , n3160, n3168);
  and g4694 (n3170, n319, n_639);
  and g4695 (n3171, n372, n_717);
  and g4699 (n3173, n426, n_744);
  and g4700 (n3174, n479, n_769);
  not g4705 (n_1927, n3176);
  and g4706 (n3177, n_182, n_1927);
  and g4707 (n3178, n319, n_692);
  and g4708 (n3179, n372, n_587);
  and g4712 (n3181, n426, n_664);
  and g4713 (n3182, n479, n_612);
  not g4718 (n_1932, n3184);
  and g4719 (n3185, \shift[6] , n_1932);
  or g4720 (\result[50] , n3177, n3185);
  and g4721 (n3187, n426, n_927);
  and g4722 (n3188, n479, n_979);
  and g4726 (n3190, n319, n_849);
  and g4727 (n3191, n372, n_954);
  not g4732 (n_1937, n3193);
  and g4733 (n3194, n_182, n_1937);
  and g4734 (n3195, n319, n_902);
  and g4735 (n3196, n426, n_797);
  and g4739 (n3198, n372, n_874);
  and g4740 (n3199, n479, n_822);
  not g4745 (n_1942, n3201);
  and g4746 (n3202, \shift[6] , n_1942);
  or g4747 (\result[51] , n3194, n3202);
  and g4748 (n3204, n426, n_1012);
  and g4749 (n3205, n319, n_999);
  and g4753 (n3207, n479, n_1024);
  and g4754 (n3208, n372, n_1029);
  not g4759 (n_1947, n3210);
  and g4760 (n3211, n_182, n_1947);
  and g4761 (n3212, n372, n_987);
  and g4762 (n3213, n479, n_992);
  and g4766 (n3215, n426, n_1004);
  and g4767 (n3216, n319, n_1017);
  not g4772 (n_1952, n3218);
  and g4773 (n3219, \shift[6] , n_1952);
  or g4774 (\result[52] , n3211, n3219);
  and g4775 (n3221, n426, n_1062);
  and g4776 (n3222, n319, n_1049);
  and g4780 (n3224, n479, n_1074);
  and g4781 (n3225, n372, n_1079);
  not g4786 (n_1957, n3227);
  and g4787 (n3228, n_182, n_1957);
  and g4788 (n3229, n372, n_1037);
  and g4789 (n3230, n479, n_1042);
  and g4793 (n3232, n426, n_1054);
  and g4794 (n3233, n319, n_1067);
  not g4799 (n_1962, n3235);
  and g4800 (n3236, \shift[6] , n_1962);
  or g4801 (\result[53] , n3228, n3236);
  and g4802 (n3238, n426, n_1112);
  and g4803 (n3239, n319, n_1099);
  and g4807 (n3241, n479, n_1124);
  and g4808 (n3242, n372, n_1129);
  not g4813 (n_1967, n3244);
  and g4814 (n3245, n_182, n_1967);
  and g4815 (n3246, n372, n_1087);
  and g4816 (n3247, n479, n_1092);
  and g4820 (n3249, n426, n_1104);
  and g4821 (n3250, n319, n_1117);
  not g4826 (n_1972, n3252);
  and g4827 (n3253, \shift[6] , n_1972);
  or g4828 (\result[54] , n3245, n3253);
  and g4829 (n3255, n426, n_1162);
  and g4830 (n3256, n372, n_1179);
  and g4834 (n3258, n319, n_1149);
  and g4835 (n3259, n479, n_1174);
  not g4840 (n_1977, n3261);
  and g4841 (n3262, n_182, n_1977);
  and g4842 (n3263, n319, n_1167);
  and g4843 (n3264, n372, n_1137);
  and g4847 (n3266, n426, n_1154);
  and g4848 (n3267, n479, n_1142);
  not g4853 (n_1982, n3269);
  and g4854 (n3270, \shift[6] , n_1982);
  or g4855 (\result[55] , n3262, n3270);
  and g4856 (n3272, n426, n_1212);
  and g4857 (n3273, n372, n_1229);
  and g4861 (n3275, n319, n_1199);
  and g4862 (n3276, n479, n_1224);
  not g4867 (n_1987, n3278);
  and g4868 (n3279, n_182, n_1987);
  and g4869 (n3280, n319, n_1217);
  and g4870 (n3281, n372, n_1187);
  and g4874 (n3283, n426, n_1204);
  and g4875 (n3284, n479, n_1192);
  not g4880 (n_1992, n3286);
  and g4881 (n3287, \shift[6] , n_1992);
  or g4882 (\result[56] , n3279, n3287);
  and g4883 (n3289, n426, n_1262);
  and g4884 (n3290, n372, n_1279);
  and g4888 (n3292, n319, n_1249);
  and g4889 (n3293, n479, n_1274);
  not g4894 (n_1997, n3295);
  and g4895 (n3296, n_182, n_1997);
  and g4896 (n3297, n319, n_1267);
  and g4897 (n3298, n372, n_1237);
  and g4901 (n3300, n426, n_1254);
  and g4902 (n3301, n479, n_1242);
  not g4907 (n_2002, n3303);
  and g4908 (n3304, \shift[6] , n_2002);
  or g4909 (\result[57] , n3296, n3304);
  and g4910 (n3306, n426, n_1312);
  and g4911 (n3307, n319, n_1299);
  and g4915 (n3309, n479, n_1324);
  and g4916 (n3310, n372, n_1329);
  not g4921 (n_2007, n3312);
  and g4922 (n3313, n_182, n_2007);
  and g4923 (n3314, n319, n_1317);
  and g4924 (n3315, n372, n_1287);
  and g4928 (n3317, n426, n_1304);
  and g4929 (n3318, n479, n_1292);
  not g4934 (n_2012, n3320);
  and g4935 (n3321, \shift[6] , n_2012);
  or g4936 (\result[58] , n3313, n3321);
  and g4937 (n3323, n426, n_1362);
  and g4938 (n3324, n319, n_1349);
  and g4942 (n3326, n479, n_1374);
  and g4943 (n3327, n372, n_1379);
  not g4948 (n_2017, n3329);
  and g4949 (n3330, n_182, n_2017);
  and g4950 (n3331, n319, n_1367);
  and g4951 (n3332, n372, n_1337);
  and g4955 (n3334, n426, n_1354);
  and g4956 (n3335, n479, n_1342);
  not g4961 (n_2022, n3337);
  and g4962 (n3338, \shift[6] , n_2022);
  or g4963 (\result[59] , n3330, n3338);
  and g4964 (n3340, n426, n_1412);
  and g4965 (n3341, n319, n_1399);
  and g4969 (n3343, n479, n_1424);
  and g4970 (n3344, n372, n_1429);
  not g4975 (n_2027, n3346);
  and g4976 (n3347, n_182, n_2027);
  and g4977 (n3348, n319, n_1417);
  and g4978 (n3349, n372, n_1387);
  and g4982 (n3351, n426, n_1404);
  and g4983 (n3352, n479, n_1392);
  not g4988 (n_2032, n3354);
  and g4989 (n3355, \shift[6] , n_2032);
  or g4990 (\result[60] , n3347, n3355);
  and g4991 (n3357, n426, n_1462);
  and g4992 (n3358, n319, n_1449);
  and g4996 (n3360, n479, n_1474);
  and g4997 (n3361, n372, n_1479);
  not g5002 (n_2037, n3363);
  and g5003 (n3364, n_182, n_2037);
  and g5004 (n3365, n319, n_1467);
  and g5005 (n3366, n372, n_1437);
  and g5009 (n3368, n426, n_1454);
  and g5010 (n3369, n479, n_1442);
  not g5015 (n_2042, n3371);
  and g5016 (n3372, \shift[6] , n_2042);
  or g5017 (\result[61] , n3364, n3372);
  and g5018 (n3374, n426, n_1512);
  and g5019 (n3375, n319, n_1499);
  and g5023 (n3377, n479, n_1524);
  and g5024 (n3378, n372, n_1529);
  not g5029 (n_2047, n3380);
  and g5030 (n3381, n_182, n_2047);
  and g5031 (n3382, n319, n_1517);
  and g5032 (n3383, n372, n_1487);
  and g5036 (n3385, n426, n_1504);
  and g5037 (n3386, n479, n_1492);
  not g5042 (n_2052, n3388);
  and g5043 (n3389, \shift[6] , n_2052);
  or g5044 (\result[62] , n3381, n3389);
  and g5045 (n3391, n426, n_1562);
  and g5046 (n3392, n319, n_1549);
  and g5050 (n3394, n479, n_1574);
  and g5051 (n3395, n372, n_1579);
  not g5056 (n_2057, n3397);
  and g5057 (n3398, n_182, n_2057);
  and g5058 (n3399, n319, n_1567);
  and g5059 (n3400, n372, n_1537);
  and g5063 (n3402, n426, n_1554);
  and g5064 (n3403, n479, n_1542);
  not g5069 (n_2062, n3405);
  and g5070 (n3406, \shift[6] , n_2062);
  or g5071 (\result[63] , n3398, n3406);
  and g5072 (n3408, n_182, n_352);
  and g5073 (n3409, \shift[6] , n_183);
  or g5074 (\result[64] , n3408, n3409);
  and g5075 (n3411, n_182, n_562);
  and g5076 (n3412, \shift[6] , n_457);
  or g5077 (\result[65] , n3411, n3412);
  and g5078 (n3414, n_182, n_772);
  and g5079 (n3415, \shift[6] , n_667);
  or g5080 (\result[66] , n3414, n3415);
  and g5081 (n3417, n_182, n_982);
  and g5082 (n3418, \shift[6] , n_877);
  or g5083 (\result[67] , n3417, n3418);
  and g5084 (n3420, n_182, n_1032);
  and g5085 (n3421, \shift[6] , n_1007);
  or g5086 (\result[68] , n3420, n3421);
  and g5087 (n3423, n_182, n_1082);
  and g5088 (n3424, \shift[6] , n_1057);
  or g5089 (\result[69] , n3423, n3424);
  and g5090 (n3426, n_182, n_1132);
  and g5091 (n3427, \shift[6] , n_1107);
  or g5092 (\result[70] , n3426, n3427);
  and g5093 (n3429, n_182, n_1182);
  and g5094 (n3430, \shift[6] , n_1157);
  or g5095 (\result[71] , n3429, n3430);
  and g5096 (n3432, n_182, n_1232);
  and g5097 (n3433, \shift[6] , n_1207);
  or g5098 (\result[72] , n3432, n3433);
  and g5099 (n3435, n_182, n_1282);
  and g5100 (n3436, \shift[6] , n_1257);
  or g5101 (\result[73] , n3435, n3436);
  and g5102 (n3438, n_182, n_1332);
  and g5103 (n3439, \shift[6] , n_1307);
  or g5104 (\result[74] , n3438, n3439);
  and g5105 (n3441, n_182, n_1382);
  and g5106 (n3442, \shift[6] , n_1357);
  or g5107 (\result[75] , n3441, n3442);
  and g5108 (n3444, n_182, n_1432);
  and g5109 (n3445, \shift[6] , n_1407);
  or g5110 (\result[76] , n3444, n3445);
  and g5111 (n3447, n_182, n_1482);
  and g5112 (n3448, \shift[6] , n_1457);
  or g5113 (\result[77] , n3447, n3448);
  and g5114 (n3450, n_182, n_1532);
  and g5115 (n3451, \shift[6] , n_1507);
  or g5116 (\result[78] , n3450, n3451);
  and g5117 (n3453, n_182, n_1582);
  and g5118 (n3454, \shift[6] , n_1557);
  or g5119 (\result[79] , n3453, n3454);
  and g5120 (n3456, n_182, n_1592);
  and g5121 (n3457, \shift[6] , n_1587);
  or g5122 (\result[80] , n3456, n3457);
  and g5123 (n3459, n_182, n_1602);
  and g5124 (n3460, \shift[6] , n_1597);
  or g5125 (\result[81] , n3459, n3460);
  and g5126 (n3462, n_182, n_1612);
  and g5127 (n3463, \shift[6] , n_1607);
  or g5128 (\result[82] , n3462, n3463);
  and g5129 (n3465, n_182, n_1622);
  and g5130 (n3466, \shift[6] , n_1617);
  or g5131 (\result[83] , n3465, n3466);
  and g5132 (n3468, n_182, n_1632);
  and g5133 (n3469, \shift[6] , n_1627);
  or g5134 (\result[84] , n3468, n3469);
  and g5135 (n3471, n_182, n_1642);
  and g5136 (n3472, \shift[6] , n_1637);
  or g5137 (\result[85] , n3471, n3472);
  and g5138 (n3474, n_182, n_1652);
  and g5139 (n3475, \shift[6] , n_1647);
  or g5140 (\result[86] , n3474, n3475);
  and g5141 (n3477, n_182, n_1662);
  and g5142 (n3478, \shift[6] , n_1657);
  or g5143 (\result[87] , n3477, n3478);
  and g5144 (n3480, n_182, n_1672);
  and g5145 (n3481, \shift[6] , n_1667);
  or g5146 (\result[88] , n3480, n3481);
  and g5147 (n3483, n_182, n_1682);
  and g5148 (n3484, \shift[6] , n_1677);
  or g5149 (\result[89] , n3483, n3484);
  and g5150 (n3486, n_182, n_1692);
  and g5151 (n3487, \shift[6] , n_1687);
  or g5152 (\result[90] , n3486, n3487);
  and g5153 (n3489, n_182, n_1702);
  and g5154 (n3490, \shift[6] , n_1697);
  or g5155 (\result[91] , n3489, n3490);
  and g5156 (n3492, n_182, n_1712);
  and g5157 (n3493, \shift[6] , n_1707);
  or g5158 (\result[92] , n3492, n3493);
  and g5159 (n3495, n_182, n_1722);
  and g5160 (n3496, \shift[6] , n_1717);
  or g5161 (\result[93] , n3495, n3496);
  and g5162 (n3498, n_182, n_1732);
  and g5163 (n3499, \shift[6] , n_1727);
  or g5164 (\result[94] , n3498, n3499);
  and g5165 (n3501, n_182, n_1742);
  and g5166 (n3502, \shift[6] , n_1737);
  or g5167 (\result[95] , n3501, n3502);
  and g5168 (n3504, n_182, n_1752);
  and g5169 (n3505, \shift[6] , n_1747);
  or g5170 (\result[96] , n3504, n3505);
  and g5171 (n3507, n_182, n_1762);
  and g5172 (n3508, \shift[6] , n_1757);
  or g5173 (\result[97] , n3507, n3508);
  and g5174 (n3510, n_182, n_1772);
  and g5175 (n3511, \shift[6] , n_1767);
  or g5176 (\result[98] , n3510, n3511);
  and g5177 (n3513, n_182, n_1782);
  and g5178 (n3514, \shift[6] , n_1777);
  or g5179 (\result[99] , n3513, n3514);
  and g5180 (n3516, n_182, n_1792);
  and g5181 (n3517, \shift[6] , n_1787);
  or g5182 (\result[100] , n3516, n3517);
  and g5183 (n3519, n_182, n_1802);
  and g5184 (n3520, \shift[6] , n_1797);
  or g5185 (\result[101] , n3519, n3520);
  and g5186 (n3522, n_182, n_1812);
  and g5187 (n3523, \shift[6] , n_1807);
  or g5188 (\result[102] , n3522, n3523);
  and g5189 (n3525, n_182, n_1822);
  and g5190 (n3526, \shift[6] , n_1817);
  or g5191 (\result[103] , n3525, n3526);
  and g5192 (n3528, n_182, n_1832);
  and g5193 (n3529, \shift[6] , n_1827);
  or g5194 (\result[104] , n3528, n3529);
  and g5195 (n3531, n_182, n_1842);
  and g5196 (n3532, \shift[6] , n_1837);
  or g5197 (\result[105] , n3531, n3532);
  and g5198 (n3534, n_182, n_1852);
  and g5199 (n3535, \shift[6] , n_1847);
  or g5200 (\result[106] , n3534, n3535);
  and g5201 (n3537, n_182, n_1862);
  and g5202 (n3538, \shift[6] , n_1857);
  or g5203 (\result[107] , n3537, n3538);
  and g5204 (n3540, n_182, n_1872);
  and g5205 (n3541, \shift[6] , n_1867);
  or g5206 (\result[108] , n3540, n3541);
  and g5207 (n3543, n_182, n_1882);
  and g5208 (n3544, \shift[6] , n_1877);
  or g5209 (\result[109] , n3543, n3544);
  and g5210 (n3546, n_182, n_1892);
  and g5211 (n3547, \shift[6] , n_1887);
  or g5212 (\result[110] , n3546, n3547);
  and g5213 (n3549, n_182, n_1902);
  and g5214 (n3550, \shift[6] , n_1897);
  or g5215 (\result[111] , n3549, n3550);
  and g5216 (n3552, n_182, n_1912);
  and g5217 (n3553, \shift[6] , n_1907);
  or g5218 (\result[112] , n3552, n3553);
  and g5219 (n3555, n_182, n_1922);
  and g5220 (n3556, \shift[6] , n_1917);
  or g5221 (\result[113] , n3555, n3556);
  and g5222 (n3558, n_182, n_1932);
  and g5223 (n3559, \shift[6] , n_1927);
  or g5224 (\result[114] , n3558, n3559);
  and g5225 (n3561, n_182, n_1942);
  and g5226 (n3562, \shift[6] , n_1937);
  or g5227 (\result[115] , n3561, n3562);
  and g5228 (n3564, n_182, n_1952);
  and g5229 (n3565, \shift[6] , n_1947);
  or g5230 (\result[116] , n3564, n3565);
  and g5231 (n3567, n_182, n_1962);
  and g5232 (n3568, \shift[6] , n_1957);
  or g5233 (\result[117] , n3567, n3568);
  and g5234 (n3570, n_182, n_1972);
  and g5235 (n3571, \shift[6] , n_1967);
  or g5236 (\result[118] , n3570, n3571);
  and g5237 (n3573, n_182, n_1982);
  and g5238 (n3574, \shift[6] , n_1977);
  or g5239 (\result[119] , n3573, n3574);
  and g5240 (n3576, n_182, n_1992);
  and g5241 (n3577, \shift[6] , n_1987);
  or g5242 (\result[120] , n3576, n3577);
  and g5243 (n3579, n_182, n_2002);
  and g5244 (n3580, \shift[6] , n_1997);
  or g5245 (\result[121] , n3579, n3580);
  and g5246 (n3582, n_182, n_2012);
  and g5247 (n3583, \shift[6] , n_2007);
  or g5248 (\result[122] , n3582, n3583);
  and g5249 (n3585, n_182, n_2022);
  and g5250 (n3586, \shift[6] , n_2017);
  or g5251 (\result[123] , n3585, n3586);
  and g5252 (n3588, n_182, n_2032);
  and g5253 (n3589, \shift[6] , n_2027);
  or g5254 (\result[124] , n3588, n3589);
  and g5255 (n3591, n_182, n_2042);
  and g5256 (n3592, \shift[6] , n_2037);
  or g5257 (\result[125] , n3591, n3592);
  and g5258 (n3594, n_182, n_2052);
  and g5259 (n3595, \shift[6] , n_2047);
  or g5260 (\result[126] , n3594, n3595);
  and g5261 (n3597, n_182, n_2062);
  and g5262 (n3598, \shift[6] , n_2057);
  or g5263 (\result[127] , n3597, n3598);
  nor g5264 (n482, n320, n373, n427, n480);
  nor g5265 (n694, n535, n587, n640, n692);
  nor g5266 (n318, n276, n289, n303, n316);
  nor g5267 (n371, n332, n344, n357, n369);
  nor g5268 (n425, n386, n398, n411, n423);
  nor g5269 (n478, n439, n451, n464, n476);
  nor g5270 (n534, n495, n507, n520, n532);
  nor g5271 (n586, n547, n559, n572, n584);
  nor g5272 (n639, n600, n612, n625, n637);
  nor g5273 (n691, n652, n664, n677, n689);
  nor g5274 (n274, n265, n267, n270, n272);
  nor g5275 (n287, n278, n280, n283, n285);
  nor g5276 (n301, n292, n294, n297, n299);
  nor g5277 (n314, n305, n307, n310, n312);
  nor g5278 (n331, n322, n324, n327, n329);
  nor g5279 (n343, n334, n336, n339, n341);
  nor g5280 (n356, n347, n349, n352, n354);
  nor g5281 (n368, n359, n361, n364, n366);
  nor g5282 (n385, n376, n378, n381, n383);
  nor g5283 (n397, n388, n390, n393, n395);
  nor g5284 (n410, n401, n403, n406, n408);
  nor g5285 (n422, n413, n415, n418, n420);
  nor g5286 (n438, n429, n431, n434, n436);
  nor g5287 (n450, n441, n443, n446, n448);
  nor g5288 (n463, n454, n456, n459, n461);
  nor g5289 (n475, n466, n468, n471, n473);
  nor g5290 (n494, n485, n487, n490, n492);
  nor g5291 (n506, n497, n499, n502, n504);
  nor g5292 (n519, n510, n512, n515, n517);
  nor g5293 (n531, n522, n524, n527, n529);
  nor g5294 (n546, n537, n539, n542, n544);
  nor g5295 (n558, n549, n551, n554, n556);
  nor g5296 (n571, n562, n564, n567, n569);
  nor g5297 (n583, n574, n576, n579, n581);
  nor g5298 (n599, n590, n592, n595, n597);
  nor g5299 (n611, n602, n604, n607, n609);
  nor g5300 (n624, n615, n617, n620, n622);
  nor g5301 (n636, n627, n629, n632, n634);
  nor g5302 (n651, n642, n644, n647, n649);
  nor g5303 (n663, n654, n656, n659, n661);
  nor g5304 (n676, n667, n669, n672, n674);
  nor g5305 (n688, n679, n681, n684, n686);
  nor g5306 (n907, n748, n800, n853, n905);
  nor g5307 (n1119, n960, n1012, n1065, n1117);
  nor g5308 (n747, n708, n720, n733, n745);
  nor g5309 (n799, n760, n772, n785, n797);
  nor g5310 (n852, n813, n825, n838, n850);
  nor g5311 (n904, n865, n877, n890, n902);
  nor g5312 (n959, n920, n932, n945, n957);
  nor g5313 (n1011, n972, n984, n997, n1009);
  nor g5314 (n1064, n1025, n1037, n1050, n1062);
  nor g5315 (n1116, n1077, n1089, n1102, n1114);
  nor g5316 (n707, n698, n700, n703, n705);
  nor g5317 (n719, n710, n712, n715, n717);
  nor g5318 (n732, n723, n725, n728, n730);
  nor g5319 (n744, n735, n737, n740, n742);
  nor g5320 (n759, n750, n752, n755, n757);
  nor g5321 (n771, n762, n764, n767, n769);
  nor g5322 (n784, n775, n777, n780, n782);
  nor g5323 (n796, n787, n789, n792, n794);
  nor g5324 (n812, n803, n805, n808, n810);
  nor g5325 (n824, n815, n817, n820, n822);
  nor g5326 (n837, n828, n830, n833, n835);
  nor g5327 (n849, n840, n842, n845, n847);
  nor g5328 (n864, n855, n857, n860, n862);
  nor g5329 (n876, n867, n869, n872, n874);
  nor g5330 (n889, n880, n882, n885, n887);
  nor g5331 (n901, n892, n894, n897, n899);
  nor g5332 (n919, n910, n912, n915, n917);
  nor g5333 (n931, n922, n924, n927, n929);
  nor g5334 (n944, n935, n937, n940, n942);
  nor g5335 (n956, n947, n949, n952, n954);
  nor g5336 (n971, n962, n964, n967, n969);
  nor g5337 (n983, n974, n976, n979, n981);
  nor g5338 (n996, n987, n989, n992, n994);
  nor g5339 (n1008, n999, n1001, n1004, n1006);
  nor g5340 (n1024, n1015, n1017, n1020, n1022);
  nor g5341 (n1036, n1027, n1029, n1032, n1034);
  nor g5342 (n1049, n1040, n1042, n1045, n1047);
  nor g5343 (n1061, n1052, n1054, n1057, n1059);
  nor g5344 (n1076, n1067, n1069, n1072, n1074);
  nor g5345 (n1088, n1079, n1081, n1084, n1086);
  nor g5346 (n1101, n1092, n1094, n1097, n1099);
  nor g5347 (n1113, n1104, n1106, n1109, n1111);
  nor g5348 (n1268, n1157, n1193, n1230, n1266);
  nor g5349 (n1416, n1305, n1341, n1378, n1414);
  nor g5350 (n1156, n1129, n1137, n1146, n1154);
  nor g5351 (n1192, n1165, n1173, n1182, n1190);
  nor g5352 (n1229, n1202, n1210, n1219, n1227);
  nor g5353 (n1265, n1238, n1246, n1255, n1263);
  nor g5354 (n1304, n1277, n1285, n1294, n1302);
  nor g5355 (n1340, n1313, n1321, n1330, n1338);
  nor g5356 (n1377, n1350, n1358, n1367, n1375);
  nor g5357 (n1413, n1386, n1394, n1403, n1411);
  nor g5358 (n1128, n1122, n1123, n1125, n1126);
  nor g5359 (n1136, n1130, n1131, n1133, n1134);
  nor g5360 (n1145, n1139, n1140, n1142, n1143);
  nor g5361 (n1153, n1147, n1148, n1150, n1151);
  nor g5362 (n1164, n1158, n1159, n1161, n1162);
  nor g5363 (n1172, n1166, n1167, n1169, n1170);
  nor g5364 (n1181, n1175, n1176, n1178, n1179);
  nor g5365 (n1189, n1183, n1184, n1186, n1187);
  nor g5366 (n1201, n1195, n1196, n1198, n1199);
  nor g5367 (n1209, n1203, n1204, n1206, n1207);
  nor g5368 (n1218, n1212, n1213, n1215, n1216);
  nor g5369 (n1226, n1220, n1221, n1223, n1224);
  nor g5370 (n1237, n1231, n1232, n1234, n1235);
  nor g5371 (n1245, n1239, n1240, n1242, n1243);
  nor g5372 (n1254, n1248, n1249, n1251, n1252);
  nor g5373 (n1262, n1256, n1257, n1259, n1260);
  nor g5374 (n1276, n1270, n1271, n1273, n1274);
  nor g5375 (n1284, n1278, n1279, n1281, n1282);
  nor g5376 (n1293, n1287, n1288, n1290, n1291);
  nor g5377 (n1301, n1295, n1296, n1298, n1299);
  nor g5378 (n1312, n1306, n1307, n1309, n1310);
  nor g5379 (n1320, n1314, n1315, n1317, n1318);
  nor g5380 (n1329, n1323, n1324, n1326, n1327);
  nor g5381 (n1337, n1331, n1332, n1334, n1335);
  nor g5382 (n1349, n1343, n1344, n1346, n1347);
  nor g5383 (n1357, n1351, n1352, n1354, n1355);
  nor g5384 (n1366, n1360, n1361, n1363, n1364);
  nor g5385 (n1374, n1368, n1369, n1371, n1372);
  nor g5386 (n1385, n1379, n1380, n1382, n1383);
  nor g5387 (n1393, n1387, n1388, n1390, n1391);
  nor g5388 (n1402, n1396, n1397, n1399, n1400);
  nor g5389 (n1410, n1404, n1405, n1407, n1408);
  nor g5390 (n1565, n1454, n1490, n1527, n1563);
  nor g5391 (n1713, n1602, n1638, n1675, n1711);
  nor g5392 (n1453, n1426, n1434, n1443, n1451);
  nor g5393 (n1489, n1462, n1470, n1479, n1487);
  nor g5394 (n1526, n1499, n1507, n1516, n1524);
  nor g5395 (n1562, n1535, n1543, n1552, n1560);
  nor g5396 (n1601, n1574, n1582, n1591, n1599);
  nor g5397 (n1637, n1610, n1618, n1627, n1635);
  nor g5398 (n1674, n1647, n1655, n1664, n1672);
  nor g5399 (n1710, n1683, n1691, n1700, n1708);
  nor g5400 (n1425, n1419, n1420, n1422, n1423);
  nor g5401 (n1433, n1427, n1428, n1430, n1431);
  nor g5402 (n1442, n1436, n1437, n1439, n1440);
  nor g5403 (n1450, n1444, n1445, n1447, n1448);
  nor g5404 (n1461, n1455, n1456, n1458, n1459);
  nor g5405 (n1469, n1463, n1464, n1466, n1467);
  nor g5406 (n1478, n1472, n1473, n1475, n1476);
  nor g5407 (n1486, n1480, n1481, n1483, n1484);
  nor g5408 (n1498, n1492, n1493, n1495, n1496);
  nor g5409 (n1506, n1500, n1501, n1503, n1504);
  nor g5410 (n1515, n1509, n1510, n1512, n1513);
  nor g5411 (n1523, n1517, n1518, n1520, n1521);
  nor g5412 (n1534, n1528, n1529, n1531, n1532);
  nor g5413 (n1542, n1536, n1537, n1539, n1540);
  nor g5414 (n1551, n1545, n1546, n1548, n1549);
  nor g5415 (n1559, n1553, n1554, n1556, n1557);
  nor g5416 (n1573, n1567, n1568, n1570, n1571);
  nor g5417 (n1581, n1575, n1576, n1578, n1579);
  nor g5418 (n1590, n1584, n1585, n1587, n1588);
  nor g5419 (n1598, n1592, n1593, n1595, n1596);
  nor g5420 (n1609, n1603, n1604, n1606, n1607);
  nor g5421 (n1617, n1611, n1612, n1614, n1615);
  nor g5422 (n1626, n1620, n1621, n1623, n1624);
  nor g5423 (n1634, n1628, n1629, n1631, n1632);
  nor g5424 (n1646, n1640, n1641, n1643, n1644);
  nor g5425 (n1654, n1648, n1649, n1651, n1652);
  nor g5426 (n1663, n1657, n1658, n1660, n1661);
  nor g5427 (n1671, n1665, n1666, n1668, n1669);
  nor g5428 (n1682, n1676, n1677, n1679, n1680);
  nor g5429 (n1690, n1684, n1685, n1687, n1688);
  nor g5430 (n1699, n1693, n1694, n1696, n1697);
  nor g5431 (n1707, n1701, n1702, n1704, n1705);
  nor g5432 (n1750, n1723, n1731, n1740, n1748);
  nor g5433 (n1786, n1759, n1767, n1776, n1784);
  nor g5434 (n1722, n1716, n1717, n1719, n1720);
  nor g5435 (n1730, n1724, n1725, n1727, n1728);
  nor g5436 (n1739, n1733, n1734, n1736, n1737);
  nor g5437 (n1747, n1741, n1742, n1744, n1745);
  nor g5438 (n1758, n1752, n1753, n1755, n1756);
  nor g5439 (n1766, n1760, n1761, n1763, n1764);
  nor g5440 (n1775, n1769, n1770, n1772, n1773);
  nor g5441 (n1783, n1777, n1778, n1780, n1781);
  nor g5442 (n1823, n1796, n1804, n1813, n1821);
  nor g5443 (n1859, n1832, n1840, n1849, n1857);
  nor g5444 (n1795, n1789, n1790, n1792, n1793);
  nor g5445 (n1803, n1797, n1798, n1800, n1801);
  nor g5446 (n1812, n1806, n1807, n1809, n1810);
  nor g5447 (n1820, n1814, n1815, n1817, n1818);
  nor g5448 (n1831, n1825, n1826, n1828, n1829);
  nor g5449 (n1839, n1833, n1834, n1836, n1837);
  nor g5450 (n1848, n1842, n1843, n1845, n1846);
  nor g5451 (n1856, n1850, n1851, n1853, n1854);
  nor g5452 (n1896, n1869, n1877, n1886, n1894);
  nor g5453 (n1932, n1905, n1913, n1922, n1930);
  nor g5454 (n1868, n1862, n1863, n1865, n1866);
  nor g5455 (n1876, n1870, n1871, n1873, n1874);
  nor g5456 (n1885, n1879, n1880, n1882, n1883);
  nor g5457 (n1893, n1887, n1888, n1890, n1891);
  nor g5458 (n1904, n1898, n1899, n1901, n1902);
  nor g5459 (n1912, n1906, n1907, n1909, n1910);
  nor g5460 (n1921, n1915, n1916, n1918, n1919);
  nor g5461 (n1929, n1923, n1924, n1926, n1927);
  nor g5462 (n1969, n1942, n1950, n1959, n1967);
  nor g5463 (n2005, n1978, n1986, n1995, n2003);
  nor g5464 (n1941, n1935, n1936, n1938, n1939);
  nor g5465 (n1949, n1943, n1944, n1946, n1947);
  nor g5466 (n1958, n1952, n1953, n1955, n1956);
  nor g5467 (n1966, n1960, n1961, n1963, n1964);
  nor g5468 (n1977, n1971, n1972, n1974, n1975);
  nor g5469 (n1985, n1979, n1980, n1982, n1983);
  nor g5470 (n1994, n1988, n1989, n1991, n1992);
  nor g5471 (n2002, n1996, n1997, n1999, n2000);
  nor g5472 (n2042, n2015, n2023, n2032, n2040);
  nor g5473 (n2078, n2051, n2059, n2068, n2076);
  nor g5474 (n2014, n2008, n2009, n2011, n2012);
  nor g5475 (n2022, n2016, n2017, n2019, n2020);
  nor g5476 (n2031, n2025, n2026, n2028, n2029);
  nor g5477 (n2039, n2033, n2034, n2036, n2037);
  nor g5478 (n2050, n2044, n2045, n2047, n2048);
  nor g5479 (n2058, n2052, n2053, n2055, n2056);
  nor g5480 (n2067, n2061, n2062, n2064, n2065);
  nor g5481 (n2075, n2069, n2070, n2072, n2073);
  nor g5482 (n2115, n2088, n2096, n2105, n2113);
  nor g5483 (n2151, n2124, n2132, n2141, n2149);
  nor g5484 (n2087, n2081, n2082, n2084, n2085);
  nor g5485 (n2095, n2089, n2090, n2092, n2093);
  nor g5486 (n2104, n2098, n2099, n2101, n2102);
  nor g5487 (n2112, n2106, n2107, n2109, n2110);
  nor g5488 (n2123, n2117, n2118, n2120, n2121);
  nor g5489 (n2131, n2125, n2126, n2128, n2129);
  nor g5490 (n2140, n2134, n2135, n2137, n2138);
  nor g5491 (n2148, n2142, n2143, n2145, n2146);
  nor g5492 (n2188, n2161, n2169, n2178, n2186);
  nor g5493 (n2224, n2197, n2205, n2214, n2222);
  nor g5494 (n2160, n2154, n2155, n2157, n2158);
  nor g5495 (n2168, n2162, n2163, n2165, n2166);
  nor g5496 (n2177, n2171, n2172, n2174, n2175);
  nor g5497 (n2185, n2179, n2180, n2182, n2183);
  nor g5498 (n2196, n2190, n2191, n2193, n2194);
  nor g5499 (n2204, n2198, n2199, n2201, n2202);
  nor g5500 (n2213, n2207, n2208, n2210, n2211);
  nor g5501 (n2221, n2215, n2216, n2218, n2219);
  nor g5502 (n2261, n2234, n2242, n2251, n2259);
  nor g5503 (n2297, n2270, n2278, n2287, n2295);
  nor g5504 (n2233, n2227, n2228, n2230, n2231);
  nor g5505 (n2241, n2235, n2236, n2238, n2239);
  nor g5506 (n2250, n2244, n2245, n2247, n2248);
  nor g5507 (n2258, n2252, n2253, n2255, n2256);
  nor g5508 (n2269, n2263, n2264, n2266, n2267);
  nor g5509 (n2277, n2271, n2272, n2274, n2275);
  nor g5510 (n2286, n2280, n2281, n2283, n2284);
  nor g5511 (n2294, n2288, n2289, n2291, n2292);
  nor g5512 (n2334, n2307, n2315, n2324, n2332);
  nor g5513 (n2370, n2343, n2351, n2360, n2368);
  nor g5514 (n2306, n2300, n2301, n2303, n2304);
  nor g5515 (n2314, n2308, n2309, n2311, n2312);
  nor g5516 (n2323, n2317, n2318, n2320, n2321);
  nor g5517 (n2331, n2325, n2326, n2328, n2329);
  nor g5518 (n2342, n2336, n2337, n2339, n2340);
  nor g5519 (n2350, n2344, n2345, n2347, n2348);
  nor g5520 (n2359, n2353, n2354, n2356, n2357);
  nor g5521 (n2367, n2361, n2362, n2364, n2365);
  nor g5522 (n2407, n2380, n2388, n2397, n2405);
  nor g5523 (n2443, n2416, n2424, n2433, n2441);
  nor g5524 (n2379, n2373, n2374, n2376, n2377);
  nor g5525 (n2387, n2381, n2382, n2384, n2385);
  nor g5526 (n2396, n2390, n2391, n2393, n2394);
  nor g5527 (n2404, n2398, n2399, n2401, n2402);
  nor g5528 (n2415, n2409, n2410, n2412, n2413);
  nor g5529 (n2423, n2417, n2418, n2420, n2421);
  nor g5530 (n2432, n2426, n2427, n2429, n2430);
  nor g5531 (n2440, n2434, n2435, n2437, n2438);
  nor g5532 (n2480, n2453, n2461, n2470, n2478);
  nor g5533 (n2516, n2489, n2497, n2506, n2514);
  nor g5534 (n2452, n2446, n2447, n2449, n2450);
  nor g5535 (n2460, n2454, n2455, n2457, n2458);
  nor g5536 (n2469, n2463, n2464, n2466, n2467);
  nor g5537 (n2477, n2471, n2472, n2474, n2475);
  nor g5538 (n2488, n2482, n2483, n2485, n2486);
  nor g5539 (n2496, n2490, n2491, n2493, n2494);
  nor g5540 (n2505, n2499, n2500, n2502, n2503);
  nor g5541 (n2513, n2507, n2508, n2510, n2511);
  nor g5542 (n2553, n2526, n2534, n2543, n2551);
  nor g5543 (n2589, n2562, n2570, n2579, n2587);
  nor g5544 (n2525, n2519, n2520, n2522, n2523);
  nor g5545 (n2533, n2527, n2528, n2530, n2531);
  nor g5546 (n2542, n2536, n2537, n2539, n2540);
  nor g5547 (n2550, n2544, n2545, n2547, n2548);
  nor g5548 (n2561, n2555, n2556, n2558, n2559);
  nor g5549 (n2569, n2563, n2564, n2566, n2567);
  nor g5550 (n2578, n2572, n2573, n2575, n2576);
  nor g5551 (n2586, n2580, n2581, n2583, n2584);
  nor g5552 (n2598, n2592, n2593, n2595, n2596);
  nor g5553 (n2606, n2600, n2601, n2603, n2604);
  nor g5554 (n2615, n2609, n2610, n2612, n2613);
  nor g5555 (n2623, n2617, n2618, n2620, n2621);
  nor g5556 (n2632, n2626, n2627, n2629, n2630);
  nor g5557 (n2640, n2634, n2635, n2637, n2638);
  nor g5558 (n2649, n2643, n2644, n2646, n2647);
  nor g5559 (n2657, n2651, n2652, n2654, n2655);
  nor g5560 (n2666, n2660, n2661, n2663, n2664);
  nor g5561 (n2674, n2668, n2669, n2671, n2672);
  nor g5562 (n2683, n2677, n2678, n2680, n2681);
  nor g5563 (n2691, n2685, n2686, n2688, n2689);
  nor g5564 (n2700, n2694, n2695, n2697, n2698);
  nor g5565 (n2708, n2702, n2703, n2705, n2706);
  nor g5566 (n2717, n2711, n2712, n2714, n2715);
  nor g5567 (n2725, n2719, n2720, n2722, n2723);
  nor g5568 (n2734, n2728, n2729, n2731, n2732);
  nor g5569 (n2742, n2736, n2737, n2739, n2740);
  nor g5570 (n2751, n2745, n2746, n2748, n2749);
  nor g5571 (n2759, n2753, n2754, n2756, n2757);
  nor g5572 (n2768, n2762, n2763, n2765, n2766);
  nor g5573 (n2776, n2770, n2771, n2773, n2774);
  nor g5574 (n2785, n2779, n2780, n2782, n2783);
  nor g5575 (n2793, n2787, n2788, n2790, n2791);
  nor g5576 (n2802, n2796, n2797, n2799, n2800);
  nor g5577 (n2810, n2804, n2805, n2807, n2808);
  nor g5578 (n2819, n2813, n2814, n2816, n2817);
  nor g5579 (n2827, n2821, n2822, n2824, n2825);
  nor g5580 (n2836, n2830, n2831, n2833, n2834);
  nor g5581 (n2844, n2838, n2839, n2841, n2842);
  nor g5582 (n2853, n2847, n2848, n2850, n2851);
  nor g5583 (n2861, n2855, n2856, n2858, n2859);
  nor g5584 (n2870, n2864, n2865, n2867, n2868);
  nor g5585 (n2878, n2872, n2873, n2875, n2876);
  nor g5586 (n2887, n2881, n2882, n2884, n2885);
  nor g5587 (n2895, n2889, n2890, n2892, n2893);
  nor g5588 (n2904, n2898, n2899, n2901, n2902);
  nor g5589 (n2912, n2906, n2907, n2909, n2910);
  nor g5590 (n2921, n2915, n2916, n2918, n2919);
  nor g5591 (n2929, n2923, n2924, n2926, n2927);
  nor g5592 (n2938, n2932, n2933, n2935, n2936);
  nor g5593 (n2946, n2940, n2941, n2943, n2944);
  nor g5594 (n2955, n2949, n2950, n2952, n2953);
  nor g5595 (n2963, n2957, n2958, n2960, n2961);
  nor g5596 (n2972, n2966, n2967, n2969, n2970);
  nor g5597 (n2980, n2974, n2975, n2977, n2978);
  nor g5598 (n2989, n2983, n2984, n2986, n2987);
  nor g5599 (n2997, n2991, n2992, n2994, n2995);
  nor g5600 (n3006, n3000, n3001, n3003, n3004);
  nor g5601 (n3014, n3008, n3009, n3011, n3012);
  nor g5602 (n3023, n3017, n3018, n3020, n3021);
  nor g5603 (n3031, n3025, n3026, n3028, n3029);
  nor g5604 (n3040, n3034, n3035, n3037, n3038);
  nor g5605 (n3048, n3042, n3043, n3045, n3046);
  nor g5606 (n3057, n3051, n3052, n3054, n3055);
  nor g5607 (n3065, n3059, n3060, n3062, n3063);
  nor g5608 (n3074, n3068, n3069, n3071, n3072);
  nor g5609 (n3082, n3076, n3077, n3079, n3080);
  nor g5610 (n3091, n3085, n3086, n3088, n3089);
  nor g5611 (n3099, n3093, n3094, n3096, n3097);
  nor g5612 (n3108, n3102, n3103, n3105, n3106);
  nor g5613 (n3116, n3110, n3111, n3113, n3114);
  nor g5614 (n3125, n3119, n3120, n3122, n3123);
  nor g5615 (n3133, n3127, n3128, n3130, n3131);
  nor g5616 (n3142, n3136, n3137, n3139, n3140);
  nor g5617 (n3150, n3144, n3145, n3147, n3148);
  nor g5618 (n3159, n3153, n3154, n3156, n3157);
  nor g5619 (n3167, n3161, n3162, n3164, n3165);
  nor g5620 (n3176, n3170, n3171, n3173, n3174);
  nor g5621 (n3184, n3178, n3179, n3181, n3182);
  nor g5622 (n3193, n3187, n3188, n3190, n3191);
  nor g5623 (n3201, n3195, n3196, n3198, n3199);
  nor g5624 (n3210, n3204, n3205, n3207, n3208);
  nor g5625 (n3218, n3212, n3213, n3215, n3216);
  nor g5626 (n3227, n3221, n3222, n3224, n3225);
  nor g5627 (n3235, n3229, n3230, n3232, n3233);
  nor g5628 (n3244, n3238, n3239, n3241, n3242);
  nor g5629 (n3252, n3246, n3247, n3249, n3250);
  nor g5630 (n3261, n3255, n3256, n3258, n3259);
  nor g5631 (n3269, n3263, n3264, n3266, n3267);
  nor g5632 (n3278, n3272, n3273, n3275, n3276);
  nor g5633 (n3286, n3280, n3281, n3283, n3284);
  nor g5634 (n3295, n3289, n3290, n3292, n3293);
  nor g5635 (n3303, n3297, n3298, n3300, n3301);
  nor g5636 (n3312, n3306, n3307, n3309, n3310);
  nor g5637 (n3320, n3314, n3315, n3317, n3318);
  nor g5638 (n3329, n3323, n3324, n3326, n3327);
  nor g5639 (n3337, n3331, n3332, n3334, n3335);
  nor g5640 (n3346, n3340, n3341, n3343, n3344);
  nor g5641 (n3354, n3348, n3349, n3351, n3352);
  nor g5642 (n3363, n3357, n3358, n3360, n3361);
  nor g5643 (n3371, n3365, n3366, n3368, n3369);
  nor g5644 (n3380, n3374, n3375, n3377, n3378);
  nor g5645 (n3388, n3382, n3383, n3385, n3386);
  nor g5646 (n3397, n3391, n3392, n3394, n3395);
  nor g5647 (n3405, n3399, n3400, n3402, n3403);
endmodule

