//# 34 inputs
//# 1 outputs
//# 32 D-type flipflops
//# 158 inverters
//# 288 gates (105 ANDs + 57 NANDs + 56 ORs + 70 NORs)

module dff (CK,Q,D);
module dff(CK,q,d);
// input CK,d;
// output reg q;
always @ (posedge CK)
q<=d;
endmodule

module s838(GND,VDD,CK,C_0,C_1,C_10,C_11,C_12,C_13,C_14,C_15,C_16,C_17,C_18,
  C_19,C_2,
  C_20,C_21,C_22,C_23,C_24,C_25,C_26,C_27,C_28,C_29,C_3,C_30,C_31,C_32,C_4,C_5,
  C_6,C_7,C_8,C_9,P_0,Z);
// input GND,VDD,CK,P_0,C_32,C_31,C_30,C_29,C_28,C_27,C_26,C_25,C_24,C_23,C_22,
  C_21,C_20,
  C_19,C_18,C_17,C_16,C_15,C_14,C_13,C_12,C_11,C_10,C_9,C_8,C_7,C_6,C_5,C_4,
  C_3,C_2,C_1,C_0;
// output Z;

  wire X_4,I12,X_3,I13,X_2,I14,X_1,I15,X_8,I110,X_7,I111,X_6,I112,X_5,I113,
    X_12,I208,X_11,I209,X_10,I210,X_9,I211,X_16,I306,X_15,I307,X_14,I308,X_13,
    I309,X_20,I404,X_19,I405,X_18,I406,X_17,I407,X_24,I502,X_23,I503,X_22,I504,
    X_21,I505,X_28,I600,X_27,I601,X_26,I602,X_25,I603,X_32,I698,X_31,I699,X_30,
    I700,X_29,I701,I73_1,I69,I73_2,I7_1,I66,I7_2,I88_1,I88_2,I48,I49,I50,I68,
    I171_1,I167,I171_2,I105_1,I164,I105_2,I186_1,I186_2,I1_2,I146,I147,I148,
    I166,I269_1,I265,I269_2,I203_1,I262,I203_2,I284_1,I284_2,I1_3,I244,I245,
    I246,I264,I367_1,I363,I367_2,I301_1,I360,I301_2,I382_1,I382_2,I1_4,I342,
    I343,I344,I362,I465_1,I461,I465_2,I399_1,I458,I399_2,I480_1,I480_2,I1_5,
    I440,I441,I442,I460,I563_1,I559,I563_2,I497_1,I556,I497_2,I578_1,I578_2,
    I1_6,I538,I539,I540,I558,I661_1,I657,I661_2,I595_1,I654,I595_2,I676_1,
    I676_2,I1_7,I636,I637,I638,I656,I693_1,I751,I693_2,I770_1,I770_2,I1_8,I736,
    I737,I749,I750,I752,I806,I807,I808,I809,I810,I819,I818,I834,I835,I836,I837,
    I838,I847,I846,I862,I863,I864,I865,I866,I875,I874,I890,I891,I892,I893,I894,
    I903,I902,I918,I919,I920,I921,I922,I931,I930,I946,I947,I948,I949,I950,I959,
    I958,I974,I975,I976,I977,I978,I987,I986,I1002,I1003,I1004,I1005,I1006,
    I1014,I1013,I1074,P_2,I1075,P_3,I1078,I1079,I1098,P_6,I1099,P_7,I1102,
    I1103,I1122,P_10,I1123,P_11,I1126,I1127,I1146,P_14,I1147,P_15,I1150,I1151,
    I1170,P_18,I1171,P_19,I1174,I1175,I1194,P_22,I1195,P_23,I1198,I1199,I1218,
    P_26,I1219,P_27,I1222,I1223,I1242,P_30,I1243,P_31,I1246,I1247,I73_3,I73_4,
    I7_3,I7_4,I88_3,I88_4,I171_3,I171_4,I105_3,I105_4,I186_3,I186_4,I269_3,
    I269_4,I203_3,I203_4,I284_3,I284_4,I367_3,I367_4,I301_3,I301_4,I382_3,
    I382_4,I465_3,I465_4,I399_3,I399_4,I480_3,I480_4,I563_3,I563_4,I497_3,
    I497_4,I578_3,I578_4,I661_3,I661_4,I595_3,I595_4,I676_3,I676_4,I693_3,
    I693_4,I770_3,I770_4,I779_1,I2_1,I2_2,I2_3,I2_4,I2_5,I2_6,I2_7,I804_2,
    I803_1,I803_2,I804_3,I803_3,I804_4,I803_4,I804_5,I803_5,I804_6,I803_6,
    I804_7,I803_7,P_5,I799_2,I800_2,I801_2,P_8,I802_2,P_9,I799_3,I800_3,I801_3,
    P_12,I802_3,P_13,I799_4,I800_4,I801_4,P_16,I802_4,P_17,I799_5,I800_5,
    I801_5,P_20,I802_5,P_21,I799_6,I800_6,I801_6,P_24,I802_6,P_25,I799_7,
    I800_7,I801_7,P_28,I802_7,P_29,I799_8,I800_8,I801_8,P_32,I802_8,I1087_1,
    P_1,I1087_2,I1111_1,I1111_2,P_4,I1135_1,I1135_2,I1159_1,I1159_2,I1183_1,
    I1183_2,I1207_1,I1207_2,I1231_1,I1231_2,I1255_1,I1255_2,I1062_9,I70_1,
    I95_1,I64,I168_1,I193_1,I162,I266_1,I291_1,I260,I364_1,I389_1,I358,I462_1,
    I487_1,I456,I560_1,I585_1,I554,I658_1,I683_1,I652,I755_1,I753,I758_1,
    I776_1,I1083_1,I1083_2,I1107_1,I1107_2,I1131_1,I1131_2,I1155_1,I1155_2,
    I1179_1,I1179_2,I1203_1,I1203_2,I1227_1,I1227_2,I1251_1,I1251_2,I1062_2,
    I1061_1,I1061_2,I1062_3,I1061_3,I1062_4,I1061_4,I1062_5,I1061_5,I1062_6,
    I1061_6,I1062_7,I1061_7,I1062_8,I1061_8,I62,I160,I258,I356,I454,I552,I650,
    I747,I816,I844,I872,I900,I928,I956,I984,I1011,I1082,I1106,I1130,I1154,
    I1178,I1202,I1226,I1250;

  dff DFF_0(CK,X_4,I12);
  dff DFF_1(CK,X_3,I13);
  dff DFF_2(CK,X_2,I14);
  dff DFF_3(CK,X_1,I15);
  dff DFF_4(CK,X_8,I110);
  dff DFF_5(CK,X_7,I111);
  dff DFF_6(CK,X_6,I112);
  dff DFF_7(CK,X_5,I113);
  dff DFF_8(CK,X_12,I208);
  dff DFF_9(CK,X_11,I209);
  dff DFF_10(CK,X_10,I210);
  dff DFF_11(CK,X_9,I211);
  dff DFF_12(CK,X_16,I306);
  dff DFF_13(CK,X_15,I307);
  dff DFF_14(CK,X_14,I308);
  dff DFF_15(CK,X_13,I309);
  dff DFF_16(CK,X_20,I404);
  dff DFF_17(CK,X_19,I405);
  dff DFF_18(CK,X_18,I406);
  dff DFF_19(CK,X_17,I407);
  dff DFF_20(CK,X_24,I502);
  dff DFF_21(CK,X_23,I503);
  dff DFF_22(CK,X_22,I504);
  dff DFF_23(CK,X_21,I505);
  dff DFF_24(CK,X_28,I600);
  dff DFF_25(CK,X_27,I601);
  dff DFF_26(CK,X_26,I602);
  dff DFF_27(CK,X_25,I603);
  dff DFF_28(CK,X_32,I698);
  dff DFF_29(CK,X_31,I699);
  dff DFF_30(CK,X_30,I700);
  dff DFF_31(CK,X_29,I701);
  not NOT_0(I73_1,I69);
  not NOT_1(I73_2,X_3);
  not NOT_2(I7_1,I66);
  not NOT_3(I7_2,X_2);
  not NOT_4(I88_1,X_1);
  not NOT_5(I88_2,P_0);
  not NOT_6(I48,P_0);
  not NOT_7(I49,X_4);
  not NOT_8(I50,X_3);
  not NOT_9(I68,I69);
  not NOT_10(I171_1,I167);
  not NOT_11(I171_2,X_7);
  not NOT_12(I105_1,I164);
  not NOT_13(I105_2,X_6);
  not NOT_14(I186_1,X_5);
  not NOT_15(I186_2,I1_2);
  not NOT_16(I146,I1_2);
  not NOT_17(I147,X_8);
  not NOT_18(I148,X_7);
  not NOT_19(I166,I167);
  not NOT_20(I269_1,I265);
  not NOT_21(I269_2,X_11);
  not NOT_22(I203_1,I262);
  not NOT_23(I203_2,X_10);
  not NOT_24(I284_1,X_9);
  not NOT_25(I284_2,I1_3);
  not NOT_26(I244,I1_3);
  not NOT_27(I245,X_12);
  not NOT_28(I246,X_11);
  not NOT_29(I264,I265);
  not NOT_30(I367_1,I363);
  not NOT_31(I367_2,X_15);
  not NOT_32(I301_1,I360);
  not NOT_33(I301_2,X_14);
  not NOT_34(I382_1,X_13);
  not NOT_35(I382_2,I1_4);
  not NOT_36(I342,I1_4);
  not NOT_37(I343,X_16);
  not NOT_38(I344,X_15);
  not NOT_39(I362,I363);
  not NOT_40(I465_1,I461);
  not NOT_41(I465_2,X_19);
  not NOT_42(I399_1,I458);
  not NOT_43(I399_2,X_18);
  not NOT_44(I480_1,X_17);
  not NOT_45(I480_2,I1_5);
  not NOT_46(I440,I1_5);
  not NOT_47(I441,X_20);
  not NOT_48(I442,X_19);
  not NOT_49(I460,I461);
  not NOT_50(I563_1,I559);
  not NOT_51(I563_2,X_23);
  not NOT_52(I497_1,I556);
  not NOT_53(I497_2,X_22);
  not NOT_54(I578_1,X_21);
  not NOT_55(I578_2,I1_6);
  not NOT_56(I538,I1_6);
  not NOT_57(I539,X_24);
  not NOT_58(I540,X_23);
  not NOT_59(I558,I559);
  not NOT_60(I661_1,I657);
  not NOT_61(I661_2,X_27);
  not NOT_62(I595_1,I654);
  not NOT_63(I595_2,X_26);
  not NOT_64(I676_1,X_25);
  not NOT_65(I676_2,I1_7);
  not NOT_66(I636,I1_7);
  not NOT_67(I637,X_28);
  not NOT_68(I638,X_27);
  not NOT_69(I656,I657);
  not NOT_70(I693_1,I751);
  not NOT_71(I693_2,X_30);
  not NOT_72(I770_1,X_29);
  not NOT_73(I770_2,I1_8);
  not NOT_74(I736,X_31);
  not NOT_75(I737,X_30);
  not NOT_76(I749,I750);
  not NOT_77(I752,I751);
  not NOT_78(I806,P_0);
  not NOT_79(I807,X_1);
  not NOT_80(I808,X_2);
  not NOT_81(I809,X_3);
  not NOT_82(I810,X_4);
  not NOT_83(I819,I818);
  not NOT_84(I834,P_0);
  not NOT_85(I835,X_5);
  not NOT_86(I836,X_6);
  not NOT_87(I837,X_7);
  not NOT_88(I838,X_8);
  not NOT_89(I847,I846);
  not NOT_90(I862,P_0);
  not NOT_91(I863,X_9);
  not NOT_92(I864,X_10);
  not NOT_93(I865,X_11);
  not NOT_94(I866,X_12);
  not NOT_95(I875,I874);
  not NOT_96(I890,P_0);
  not NOT_97(I891,X_13);
  not NOT_98(I892,X_14);
  not NOT_99(I893,X_15);
  not NOT_100(I894,X_16);
  not NOT_101(I903,I902);
  not NOT_102(I918,P_0);
  not NOT_103(I919,X_17);
  not NOT_104(I920,X_18);
  not NOT_105(I921,X_19);
  not NOT_106(I922,X_20);
  not NOT_107(I931,I930);
  not NOT_108(I946,P_0);
  not NOT_109(I947,X_21);
  not NOT_110(I948,X_22);
  not NOT_111(I949,X_23);
  not NOT_112(I950,X_24);
  not NOT_113(I959,I958);
  not NOT_114(I974,P_0);
  not NOT_115(I975,X_25);
  not NOT_116(I976,X_26);
  not NOT_117(I977,X_27);
  not NOT_118(I978,X_28);
  not NOT_119(I987,I986);
  not NOT_120(I1002,P_0);
  not NOT_121(I1003,X_29);
  not NOT_122(I1004,X_30);
  not NOT_123(I1005,X_31);
  not NOT_124(I1006,X_32);
  not NOT_125(I1014,I1013);
  not NOT_126(I1074,P_2);
  not NOT_127(I1075,P_3);
  not NOT_128(I1078,C_2);
  not NOT_129(I1079,C_3);
  not NOT_130(I1098,P_6);
  not NOT_131(I1099,P_7);
  not NOT_132(I1102,C_6);
  not NOT_133(I1103,C_7);
  not NOT_134(I1122,P_10);
  not NOT_135(I1123,P_11);
  not NOT_136(I1126,C_10);
  not NOT_137(I1127,C_11);
  not NOT_138(I1146,P_14);
  not NOT_139(I1147,P_15);
  not NOT_140(I1150,C_14);
  not NOT_141(I1151,C_15);
  not NOT_142(I1170,P_18);
  not NOT_143(I1171,P_19);
  not NOT_144(I1174,C_18);
  not NOT_145(I1175,C_19);
  not NOT_146(I1194,P_22);
  not NOT_147(I1195,P_23);
  not NOT_148(I1198,C_22);
  not NOT_149(I1199,C_23);
  not NOT_150(I1218,P_26);
  not NOT_151(I1219,P_27);
  not NOT_152(I1222,C_26);
  not NOT_153(I1223,C_27);
  not NOT_154(I1242,P_30);
  not NOT_155(I1243,P_31);
  not NOT_156(I1246,C_30);
  not NOT_157(I1247,C_31);
  and AND2_0(I73_3,I69,I73_2);
  and AND2_1(I73_4,X_3,I73_1);
  and AND2_2(I7_3,I66,I7_2);
  and AND2_3(I7_4,X_2,I7_1);
  and AND2_4(I88_3,X_1,I88_2);
  and AND2_5(I88_4,P_0,I88_1);
  and AND2_6(I171_3,I167,I171_2);
  and AND2_7(I171_4,X_7,I171_1);
  and AND2_8(I105_3,I164,I105_2);
  and AND2_9(I105_4,X_6,I105_1);
  and AND2_10(I186_3,X_5,I186_2);
  and AND2_11(I186_4,I1_2,I186_1);
  and AND2_12(I269_3,I265,I269_2);
  and AND2_13(I269_4,X_11,I269_1);
  and AND2_14(I203_3,I262,I203_2);
  and AND2_15(I203_4,X_10,I203_1);
  and AND2_16(I284_3,X_9,I284_2);
  and AND2_17(I284_4,I1_3,I284_1);
  and AND2_18(I367_3,I363,I367_2);
  and AND2_19(I367_4,X_15,I367_1);
  and AND2_20(I301_3,I360,I301_2);
  and AND2_21(I301_4,X_14,I301_1);
  and AND2_22(I382_3,X_13,I382_2);
  and AND2_23(I382_4,I1_4,I382_1);
  and AND2_24(I465_3,I461,I465_2);
  and AND2_25(I465_4,X_19,I465_1);
  and AND2_26(I399_3,I458,I399_2);
  and AND2_27(I399_4,X_18,I399_1);
  and AND2_28(I480_3,X_17,I480_2);
  and AND2_29(I480_4,I1_5,I480_1);
  and AND2_30(I563_3,I559,I563_2);
  and AND2_31(I563_4,X_23,I563_1);
  and AND2_32(I497_3,I556,I497_2);
  and AND2_33(I497_4,X_22,I497_1);
  and AND2_34(I578_3,X_21,I578_2);
  and AND2_35(I578_4,I1_6,I578_1);
  and AND2_36(I661_3,I657,I661_2);
  and AND2_37(I661_4,X_27,I661_1);
  and AND2_38(I595_3,I654,I595_2);
  and AND2_39(I595_4,X_26,I595_1);
  and AND2_40(I676_3,X_25,I676_2);
  and AND2_41(I676_4,I1_7,I676_1);
  and AND2_42(I693_3,I751,I693_2);
  and AND2_43(I693_4,X_30,I693_1);
  and AND2_44(I770_3,X_29,I770_2);
  and AND2_45(I770_4,I1_8,I770_1);
  and AND2_46(I779_1,I752,X_30);
  and AND2_47(I1_2,I2_1,P_0);
  and AND2_48(I1_3,I2_2,I1_2);
  and AND2_49(I1_4,I2_3,I1_3);
  and AND2_50(I1_5,I2_4,I1_4);
  and AND2_51(I1_6,I2_5,I1_5);
  and AND2_52(I1_7,I2_6,I1_6);
  and AND2_53(I1_8,I2_7,I1_7);
  and AND2_54(I804_2,I803_1,I803_2);
  and AND2_55(I804_3,I804_2,I803_3);
  and AND2_56(I804_4,I804_3,I803_4);
  and AND2_57(I804_5,I804_4,I803_5);
  and AND2_58(I804_6,I804_5,I803_6);
  and AND2_59(I804_7,I804_6,I803_7);
  and AND2_60(P_5,I803_1,I799_2);
  and AND2_61(P_6,I803_1,I800_2);
  and AND2_62(P_7,I803_1,I801_2);
  and AND2_63(P_8,I803_1,I802_2);
  and AND2_64(P_9,I804_2,I799_3);
  and AND2_65(P_10,I804_2,I800_3);
  and AND2_66(P_11,I804_2,I801_3);
  and AND2_67(P_12,I804_2,I802_3);
  and AND2_68(P_13,I804_3,I799_4);
  and AND2_69(P_14,I804_3,I800_4);
  and AND2_70(P_15,I804_3,I801_4);
  and AND2_71(P_16,I804_3,I802_4);
  and AND2_72(P_17,I804_4,I799_5);
  and AND2_73(P_18,I804_4,I800_5);
  and AND2_74(P_19,I804_4,I801_5);
  and AND2_75(P_20,I804_4,I802_5);
  and AND2_76(P_21,I804_5,I799_6);
  and AND2_77(P_22,I804_5,I800_6);
  and AND2_78(P_23,I804_5,I801_6);
  and AND2_79(P_24,I804_5,I802_6);
  and AND2_80(P_25,I804_6,I799_7);
  and AND2_81(P_26,I804_6,I800_7);
  and AND2_82(P_27,I804_6,I801_7);
  and AND2_83(P_28,I804_6,I802_7);
  and AND2_84(P_29,I804_7,I799_8);
  and AND2_85(P_30,I804_7,I800_8);
  and AND2_86(P_31,I804_7,I801_8);
  and AND2_87(P_32,I804_7,I802_8);
  and AND2_88(I1087_1,P_1,C_1);
  and AND2_89(I1087_2,P_0,C_0);
  and AND2_90(I1111_1,P_5,C_5);
  and AND2_91(I1111_2,P_4,C_4);
  and AND2_92(I1135_1,P_9,C_9);
  and AND2_93(I1135_2,P_8,C_8);
  and AND2_94(I1159_1,P_13,C_13);
  and AND2_95(I1159_2,P_12,C_12);
  and AND2_96(I1183_1,P_17,C_17);
  and AND2_97(I1183_2,P_16,C_16);
  and AND2_98(I1207_1,P_21,C_21);
  and AND2_99(I1207_2,P_20,C_20);
  and AND2_100(I1231_1,P_25,C_25);
  and AND2_101(I1231_2,P_24,C_24);
  and AND2_102(I1255_1,P_29,C_29);
  and AND2_103(I1255_2,P_28,C_28);
  and AND2_104(I1062_9,P_32,C_32);
  or OR3_0(I70_1,I68,X_4,I50);
  or OR2_0(I13,I73_3,I73_4);
  or OR2_1(I15,I88_3,I88_4);
  or OR3_1(I95_1,I64,I50,I48);
  or OR3_2(I168_1,I166,X_8,I148);
  or OR2_2(I111,I171_3,I171_4);
  or OR2_3(I113,I186_3,I186_4);
  or OR3_3(I193_1,I162,I148,I146);
  or OR3_4(I266_1,I264,X_12,I246);
  or OR2_4(I209,I269_3,I269_4);
  or OR2_5(I211,I284_3,I284_4);
  or OR3_5(I291_1,I260,I246,I244);
  or OR3_6(I364_1,I362,X_16,I344);
  or OR2_6(I307,I367_3,I367_4);
  or OR2_7(I309,I382_3,I382_4);
  or OR3_7(I389_1,I358,I344,I342);
  or OR3_8(I462_1,I460,X_20,I442);
  or OR2_8(I405,I465_3,I465_4);
  or OR2_9(I407,I480_3,I480_4);
  or OR3_9(I487_1,I456,I442,I440);
  or OR3_10(I560_1,I558,X_24,I540);
  or OR2_10(I503,I563_3,I563_4);
  or OR2_11(I505,I578_3,I578_4);
  or OR3_11(I585_1,I554,I540,I538);
  or OR3_12(I658_1,I656,X_28,I638);
  or OR2_12(I601,I661_3,I661_4);
  or OR2_13(I603,I676_3,I676_4);
  or OR3_13(I683_1,I652,I638,I636);
  or OR3_14(I755_1,I753,X_32,I736);
  or OR2_14(I758_1,I753,X_31);
  or OR2_15(I701,I770_3,I770_4);
  or OR3_15(I776_1,I751,I737,I736);
  or OR2_16(I1083_1,I1075,I1079);
  or OR2_17(I1083_2,I1074,I1078);
  or OR2_18(I1107_1,I1099,I1103);
  or OR2_19(I1107_2,I1098,I1102);
  or OR2_20(I1131_1,I1123,I1127);
  or OR2_21(I1131_2,I1122,I1126);
  or OR2_22(I1155_1,I1147,I1151);
  or OR2_23(I1155_2,I1146,I1150);
  or OR2_24(I1179_1,I1171,I1175);
  or OR2_25(I1179_2,I1170,I1174);
  or OR2_26(I1203_1,I1195,I1199);
  or OR2_27(I1203_2,I1194,I1198);
  or OR2_28(I1227_1,I1219,I1223);
  or OR2_29(I1227_2,I1218,I1222);
  or OR2_30(I1251_1,I1243,I1247);
  or OR2_31(I1251_2,I1242,I1246);
  or OR2_32(I1062_2,I1061_1,I1061_2);
  or OR2_33(I1062_3,I1062_2,I1061_3);
  or OR2_34(I1062_4,I1062_3,I1061_4);
  or OR2_35(I1062_5,I1062_4,I1061_5);
  or OR2_36(I1062_6,I1062_5,I1061_6);
  or OR2_37(I1062_7,I1062_6,I1061_7);
  or OR2_38(I1062_8,I1062_7,I1061_8);
  or OR2_39(Z,I1062_8,I1062_9);
  nand NAND2_0(I12,I70_1,I62);
  nand NAND2_1(I62,I95_1,X_4);
  nand NAND2_2(I64,X_1,X_2);
  nand NAND2_3(I66,X_1,P_0);
  nand NAND2_4(I110,I168_1,I160);
  nand NAND2_5(I160,I193_1,X_8);
  nand NAND2_6(I162,X_5,X_6);
  nand NAND2_7(I164,X_5,I1_2);
  nand NAND2_8(I208,I266_1,I258);
  nand NAND2_9(I258,I291_1,X_12);
  nand NAND2_10(I260,X_9,X_10);
  nand NAND2_11(I262,X_9,I1_3);
  nand NAND2_12(I306,I364_1,I356);
  nand NAND2_13(I356,I389_1,X_16);
  nand NAND2_14(I358,X_13,X_14);
  nand NAND2_15(I360,X_13,I1_4);
  nand NAND2_16(I404,I462_1,I454);
  nand NAND2_17(I454,I487_1,X_20);
  nand NAND2_18(I456,X_17,X_18);
  nand NAND2_19(I458,X_17,I1_5);
  nand NAND2_20(I502,I560_1,I552);
  nand NAND2_21(I552,I585_1,X_24);
  nand NAND2_22(I554,X_21,X_22);
  nand NAND2_23(I556,X_21,I1_6);
  nand NAND2_24(I600,I658_1,I650);
  nand NAND2_25(I650,I683_1,X_28);
  nand NAND2_26(I652,X_25,X_26);
  nand NAND2_27(I654,X_25,I1_7);
  nand NAND2_28(I698,I755_1,I747);
  nand NAND2_29(I699,I758_1,I749);
  nand NAND2_30(I747,I776_1,X_32);
  nand NAND2_31(I751,X_29,I1_8);
  nand NAND2_32(I753,I752,X_30);
  nand NAND2_33(I816,I819,I808);
  nand NAND2_34(I818,I807,P_0);
  nand NAND2_35(I844,I847,I836);
  nand NAND2_36(I846,I835,P_0);
  nand NAND2_37(I872,I875,I864);
  nand NAND2_38(I874,I863,P_0);
  nand NAND2_39(I900,I903,I892);
  nand NAND2_40(I902,I891,P_0);
  nand NAND2_41(I928,I931,I920);
  nand NAND2_42(I930,I919,P_0);
  nand NAND2_43(I956,I959,I948);
  nand NAND2_44(I958,I947,P_0);
  nand NAND2_45(I984,I987,I976);
  nand NAND2_46(I986,I975,P_0);
  nand NAND2_47(I1011,I1014,I1004);
  nand NAND2_48(I1013,I1003,P_0);
  nand NAND3_0(I1061_1,I1083_1,I1083_2,I1082);
  nand NAND3_1(I1061_2,I1107_1,I1107_2,I1106);
  nand NAND3_2(I1061_3,I1131_1,I1131_2,I1130);
  nand NAND3_3(I1061_4,I1155_1,I1155_2,I1154);
  nand NAND3_4(I1061_5,I1179_1,I1179_2,I1178);
  nand NAND3_5(I1061_6,I1203_1,I1203_2,I1202);
  nand NAND3_6(I1061_7,I1227_1,I1227_2,I1226);
  nand NAND3_7(I1061_8,I1251_1,I1251_2,I1250);
  nor NOR2_0(I14,I7_3,I7_4);
  nor NOR3_0(I2_1,I64,I49,I50);
  nor NOR2_1(I69,I64,I48);
  nor NOR2_2(I112,I105_3,I105_4);
  nor NOR3_1(I2_2,I162,I147,I148);
  nor NOR2_3(I167,I162,I146);
  nor NOR2_4(I210,I203_3,I203_4);
  nor NOR3_2(I2_3,I260,I245,I246);
  nor NOR2_5(I265,I260,I244);
  nor NOR2_6(I308,I301_3,I301_4);
  nor NOR3_3(I2_4,I358,I343,I344);
  nor NOR2_7(I363,I358,I342);
  nor NOR2_8(I406,I399_3,I399_4);
  nor NOR3_4(I2_5,I456,I441,I442);
  nor NOR2_9(I461,I456,I440);
  nor NOR2_10(I504,I497_3,I497_4);
  nor NOR3_5(I2_6,I554,I539,I540);
  nor NOR2_11(I559,I554,I538);
  nor NOR2_12(I602,I595_3,I595_4);
  nor NOR3_6(I2_7,I652,I637,I638);
  nor NOR2_13(I657,I652,I636);
  nor NOR2_14(I700,I693_3,I693_4);
  nor NOR2_15(I750,I736,I779_1);
  nor NOR2_16(P_1,I806,I807);
  nor NOR2_17(P_2,I808,I818);
  nor NOR2_18(P_3,I809,I816);
  nor NOR3_7(P_4,X_3,I816,I810);
  nor NOR4_0(I803_1,X_4,X_2,X_3,X_1);
  nor NOR2_19(I799_2,I834,I835);
  nor NOR2_20(I800_2,I836,I846);
  nor NOR2_21(I801_2,I837,I844);
  nor NOR3_8(I802_2,X_7,I844,I838);
  nor NOR4_1(I803_2,X_8,X_6,X_7,X_5);
  nor NOR2_22(I799_3,I862,I863);
  nor NOR2_23(I800_3,I864,I874);
  nor NOR2_24(I801_3,I865,I872);
  nor NOR3_9(I802_3,X_11,I872,I866);
  nor NOR4_2(I803_3,X_12,X_10,X_11,X_9);
  nor NOR2_25(I799_4,I890,I891);
  nor NOR2_26(I800_4,I892,I902);
  nor NOR2_27(I801_4,I893,I900);
  nor NOR3_10(I802_4,X_15,I900,I894);
  nor NOR4_3(I803_4,X_16,X_14,X_15,X_13);
  nor NOR2_28(I799_5,I918,I919);
  nor NOR2_29(I800_5,I920,I930);
  nor NOR2_30(I801_5,I921,I928);
  nor NOR3_11(I802_5,X_19,I928,I922);
  nor NOR4_4(I803_5,X_20,X_18,X_19,X_17);
  nor NOR2_31(I799_6,I946,I947);
  nor NOR2_32(I800_6,I948,I958);
  nor NOR2_33(I801_6,I949,I956);
  nor NOR3_12(I802_6,X_23,I956,I950);
  nor NOR4_5(I803_6,X_24,X_22,X_23,X_21);
  nor NOR2_34(I799_7,I974,I975);
  nor NOR2_35(I800_7,I976,I986);
  nor NOR2_36(I801_7,I977,I984);
  nor NOR3_13(I802_7,X_27,I984,I978);
  nor NOR4_6(I803_7,X_28,X_26,X_27,X_25);
  nor NOR2_37(I799_8,I1002,I1003);
  nor NOR2_38(I800_8,I1004,I1013);
  nor NOR2_39(I801_8,I1005,I1011);
  nor NOR3_14(I802_8,X_31,I1011,I1006);
  nor NOR2_40(I1082,I1087_1,I1087_2);
  nor NOR2_41(I1106,I1111_1,I1111_2);
  nor NOR2_42(I1130,I1135_1,I1135_2);
  nor NOR2_43(I1154,I1159_1,I1159_2);
  nor NOR2_44(I1178,I1183_1,I1183_2);
  nor NOR2_45(I1202,I1207_1,I1207_2);
  nor NOR2_46(I1226,I1231_1,I1231_2);
  nor NOR2_47(I1250,I1255_1,I1255_2);

endmodule

