
module arbiter(\priority[0] , \priority[1] , \priority[2] ,
     \priority[3] , \priority[4] , \priority[5] , \priority[6] ,
     \priority[7] , \priority[8] , \priority[9] , \priority[10] ,
     \priority[11] , \priority[12] , \priority[13] , \priority[14] ,
     \priority[15] , \priority[16] , \priority[17] , \priority[18] ,
     \priority[19] , \priority[20] , \priority[21] , \priority[22] ,
     \priority[23] , \priority[24] , \priority[25] , \priority[26] ,
     \priority[27] , \priority[28] , \priority[29] , \priority[30] ,
     \priority[31] , \priority[32] , \priority[33] , \priority[34] ,
     \priority[35] , \priority[36] , \priority[37] , \priority[38] ,
     \priority[39] , \priority[40] , \priority[41] , \priority[42] ,
     \priority[43] , \priority[44] , \priority[45] , \priority[46] ,
     \priority[47] , \priority[48] , \priority[49] , \priority[50] ,
     \priority[51] , \priority[52] , \priority[53] , \priority[54] ,
     \priority[55] , \priority[56] , \priority[57] , \priority[58] ,
     \priority[59] , \priority[60] , \priority[61] , \priority[62] ,
     \priority[63] , \priority[64] , \priority[65] , \priority[66] ,
     \priority[67] , \priority[68] , \priority[69] , \priority[70] ,
     \priority[71] , \priority[72] , \priority[73] , \priority[74] ,
     \priority[75] , \priority[76] , \priority[77] , \priority[78] ,
     \priority[79] , \priority[80] , \priority[81] , \priority[82] ,
     \priority[83] , \priority[84] , \priority[85] , \priority[86] ,
     \priority[87] , \priority[88] , \priority[89] , \priority[90] ,
     \priority[91] , \priority[92] , \priority[93] , \priority[94] ,
     \priority[95] , \priority[96] , \priority[97] , \priority[98] ,
     \priority[99] , \priority[100] , \priority[101] , \priority[102] ,
     \priority[103] , \priority[104] , \priority[105] , \priority[106]
     , \priority[107] , \priority[108] , \priority[109] ,
     \priority[110] , \priority[111] , \priority[112] , \priority[113]
     , \priority[114] , \priority[115] , \priority[116] ,
     \priority[117] , \priority[118] , \priority[119] , \priority[120]
     , \priority[121] , \priority[122] , \priority[123] ,
     \priority[124] , \priority[125] , \priority[126] , \priority[127]
     , \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] ,
     \req[6] , \req[7] , \req[8] , \req[9] , \req[10] , \req[11] ,
     \req[12] , \req[13] , \req[14] , \req[15] , \req[16] , \req[17] ,
     \req[18] , \req[19] , \req[20] , \req[21] , \req[22] , \req[23] ,
     \req[24] , \req[25] , \req[26] , \req[27] , \req[28] , \req[29] ,
     \req[30] , \req[31] , \req[32] , \req[33] , \req[34] , \req[35] ,
     \req[36] , \req[37] , \req[38] , \req[39] , \req[40] , \req[41] ,
     \req[42] , \req[43] , \req[44] , \req[45] , \req[46] , \req[47] ,
     \req[48] , \req[49] , \req[50] , \req[51] , \req[52] , \req[53] ,
     \req[54] , \req[55] , \req[56] , \req[57] , \req[58] , \req[59] ,
     \req[60] , \req[61] , \req[62] , \req[63] , \req[64] , \req[65] ,
     \req[66] , \req[67] , \req[68] , \req[69] , \req[70] , \req[71] ,
     \req[72] , \req[73] , \req[74] , \req[75] , \req[76] , \req[77] ,
     \req[78] , \req[79] , \req[80] , \req[81] , \req[82] , \req[83] ,
     \req[84] , \req[85] , \req[86] , \req[87] , \req[88] , \req[89] ,
     \req[90] , \req[91] , \req[92] , \req[93] , \req[94] , \req[95] ,
     \req[96] , \req[97] , \req[98] , \req[99] , \req[100] , \req[101]
     , \req[102] , \req[103] , \req[104] , \req[105] , \req[106] ,
     \req[107] , \req[108] , \req[109] , \req[110] , \req[111] ,
     \req[112] , \req[113] , \req[114] , \req[115] , \req[116] ,
     \req[117] , \req[118] , \req[119] , \req[120] , \req[121] ,
     \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
     \req[127] , \grant[0] , \grant[1] , \grant[2] , \grant[3] ,
     \grant[4] , \grant[5] , \grant[6] , \grant[7] , \grant[8] ,
     \grant[9] , \grant[10] , \grant[11] , \grant[12] , \grant[13] ,
     \grant[14] , \grant[15] , \grant[16] , \grant[17] , \grant[18] ,
     \grant[19] , \grant[20] , \grant[21] , \grant[22] , \grant[23] ,
     \grant[24] , \grant[25] , \grant[26] , \grant[27] , \grant[28] ,
     \grant[29] , \grant[30] , \grant[31] , \grant[32] , \grant[33] ,
     \grant[34] , \grant[35] , \grant[36] , \grant[37] , \grant[38] ,
     \grant[39] , \grant[40] , \grant[41] , \grant[42] , \grant[43] ,
     \grant[44] , \grant[45] , \grant[46] , \grant[47] , \grant[48] ,
     \grant[49] , \grant[50] , \grant[51] , \grant[52] , \grant[53] ,
     \grant[54] , \grant[55] , \grant[56] , \grant[57] , \grant[58] ,
     \grant[59] , \grant[60] , \grant[61] , \grant[62] , \grant[63] ,
     \grant[64] , \grant[65] , \grant[66] , \grant[67] , \grant[68] ,
     \grant[69] , \grant[70] , \grant[71] , \grant[72] , \grant[73] ,
     \grant[74] , \grant[75] , \grant[76] , \grant[77] , \grant[78] ,
     \grant[79] , \grant[80] , \grant[81] , \grant[82] , \grant[83] ,
     \grant[84] , \grant[85] , \grant[86] , \grant[87] , \grant[88] ,
     \grant[89] , \grant[90] , \grant[91] , \grant[92] , \grant[93] ,
     \grant[94] , \grant[95] , \grant[96] , \grant[97] , \grant[98] ,
     \grant[99] , \grant[100] , \grant[101] , \grant[102] , \grant[103]
     , \grant[104] , \grant[105] , \grant[106] , \grant[107] ,
     \grant[108] , \grant[109] , \grant[110] , \grant[111] ,
     \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
     \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
     \grant[120] , \grant[121] , \grant[122] , \grant[123] ,
     \grant[124] , \grant[125] , \grant[126] , \grant[127] , anyGrant);
  input \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
       \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
       \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
       \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
       \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
       \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
       \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
       \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
       \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
       \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
       \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
       \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
       \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
       \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
       \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
       \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
       \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
       \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
       \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
       \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
       \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
       \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
       \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
       \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
       \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
       \priority[100] , \priority[101] , \priority[102] ,
       \priority[103] , \priority[104] , \priority[105] ,
       \priority[106] , \priority[107] , \priority[108] ,
       \priority[109] , \priority[110] , \priority[111] ,
       \priority[112] , \priority[113] , \priority[114] ,
       \priority[115] , \priority[116] , \priority[117] ,
       \priority[118] , \priority[119] , \priority[120] ,
       \priority[121] , \priority[122] , \priority[123] ,
       \priority[124] , \priority[125] , \priority[126] ,
       \priority[127] , \req[0] , \req[1] , \req[2] , \req[3] , \req[4]
       , \req[5] , \req[6] , \req[7] , \req[8] , \req[9] , \req[10] ,
       \req[11] , \req[12] , \req[13] , \req[14] , \req[15] , \req[16]
       , \req[17] , \req[18] , \req[19] , \req[20] , \req[21] ,
       \req[22] , \req[23] , \req[24] , \req[25] , \req[26] , \req[27]
       , \req[28] , \req[29] , \req[30] , \req[31] , \req[32] ,
       \req[33] , \req[34] , \req[35] , \req[36] , \req[37] , \req[38]
       , \req[39] , \req[40] , \req[41] , \req[42] , \req[43] ,
       \req[44] , \req[45] , \req[46] , \req[47] , \req[48] , \req[49]
       , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
       \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60]
       , \req[61] , \req[62] , \req[63] , \req[64] , \req[65] ,
       \req[66] , \req[67] , \req[68] , \req[69] , \req[70] , \req[71]
       , \req[72] , \req[73] , \req[74] , \req[75] , \req[76] ,
       \req[77] , \req[78] , \req[79] , \req[80] , \req[81] , \req[82]
       , \req[83] , \req[84] , \req[85] , \req[86] , \req[87] ,
       \req[88] , \req[89] , \req[90] , \req[91] , \req[92] , \req[93]
       , \req[94] , \req[95] , \req[96] , \req[97] , \req[98] ,
       \req[99] , \req[100] , \req[101] , \req[102] , \req[103] ,
       \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
       \req[109] , \req[110] , \req[111] , \req[112] , \req[113] ,
       \req[114] , \req[115] , \req[116] , \req[117] , \req[118] ,
       \req[119] , \req[120] , \req[121] , \req[122] , \req[123] ,
       \req[124] , \req[125] , \req[126] , \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
       \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
       \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
       \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
       \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
       \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
       \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
       \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
       \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
       \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
       \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
       \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
       \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
       \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
       \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
       \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
       \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
       \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
       \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
       \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
       \grant[100] , \grant[101] , \grant[102] , \grant[103] ,
       \grant[104] , \grant[105] , \grant[106] , \grant[107] ,
       \grant[108] , \grant[109] , \grant[110] , \grant[111] ,
       \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
       \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
       \grant[120] , \grant[121] , \grant[122] , \grant[123] ,
       \grant[124] , \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
       \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
       \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
       \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
       \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
       \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
       \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
       \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
       \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
       \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
       \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
       \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
       \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
       \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
       \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
       \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
       \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
       \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
       \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
       \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
       \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
       \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
       \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
       \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
       \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
       \priority[100] , \priority[101] , \priority[102] ,
       \priority[103] , \priority[104] , \priority[105] ,
       \priority[106] , \priority[107] , \priority[108] ,
       \priority[109] , \priority[110] , \priority[111] ,
       \priority[112] , \priority[113] , \priority[114] ,
       \priority[115] , \priority[116] , \priority[117] ,
       \priority[118] , \priority[119] , \priority[120] ,
       \priority[121] , \priority[122] , \priority[123] ,
       \priority[124] , \priority[125] , \priority[126] ,
       \priority[127] , \req[0] , \req[1] , \req[2] , \req[3] , \req[4]
       , \req[5] , \req[6] , \req[7] , \req[8] , \req[9] , \req[10] ,
       \req[11] , \req[12] , \req[13] , \req[14] , \req[15] , \req[16]
       , \req[17] , \req[18] , \req[19] , \req[20] , \req[21] ,
       \req[22] , \req[23] , \req[24] , \req[25] , \req[26] , \req[27]
       , \req[28] , \req[29] , \req[30] , \req[31] , \req[32] ,
       \req[33] , \req[34] , \req[35] , \req[36] , \req[37] , \req[38]
       , \req[39] , \req[40] , \req[41] , \req[42] , \req[43] ,
       \req[44] , \req[45] , \req[46] , \req[47] , \req[48] , \req[49]
       , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
       \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60]
       , \req[61] , \req[62] , \req[63] , \req[64] , \req[65] ,
       \req[66] , \req[67] , \req[68] , \req[69] , \req[70] , \req[71]
       , \req[72] , \req[73] , \req[74] , \req[75] , \req[76] ,
       \req[77] , \req[78] , \req[79] , \req[80] , \req[81] , \req[82]
       , \req[83] , \req[84] , \req[85] , \req[86] , \req[87] ,
       \req[88] , \req[89] , \req[90] , \req[91] , \req[92] , \req[93]
       , \req[94] , \req[95] , \req[96] , \req[97] , \req[98] ,
       \req[99] , \req[100] , \req[101] , \req[102] , \req[103] ,
       \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
       \req[109] , \req[110] , \req[111] , \req[112] , \req[113] ,
       \req[114] , \req[115] , \req[116] , \req[117] , \req[118] ,
       \req[119] , \req[120] , \req[121] , \req[122] , \req[123] ,
       \req[124] , \req[125] , \req[126] , \req[127] ;
  wire \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
       \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
       \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
       \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
       \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
       \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
       \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
       \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
       \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
       \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
       \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
       \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
       \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
       \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
       \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
       \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
       \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
       \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
       \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
       \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
       \grant[100] , \grant[101] , \grant[102] , \grant[103] ,
       \grant[104] , \grant[105] , \grant[106] , \grant[107] ,
       \grant[108] , \grant[109] , \grant[110] , \grant[111] ,
       \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
       \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
       \grant[120] , \grant[121] , \grant[122] , \grant[123] ,
       \grant[124] , \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire n386, n387, n388, n389, n390, n391, n392, n393;
  wire n394, n395, n396, n397, n398, n399, n400, n401;
  wire n402, n403, n404, n405, n406, n407, n408, n409;
  wire n410, n411, n412, n413, n414, n415, n416, n417;
  wire n418, n419, n420, n421, n422, n423, n424, n425;
  wire n426, n427, n428, n429, n430, n431, n432, n433;
  wire n434, n435, n436, n437, n438, n439, n440, n441;
  wire n442, n443, n444, n445, n446, n447, n448, n449;
  wire n450, n451, n452, n453, n454, n455, n456, n457;
  wire n458, n459, n460, n461, n462, n463, n464, n465;
  wire n466, n467, n468, n469, n470, n471, n472, n473;
  wire n474, n475, n476, n477, n478, n479, n480, n481;
  wire n482, n483, n484, n485, n486, n487, n488, n489;
  wire n490, n491, n492, n493, n494, n495, n496, n497;
  wire n498, n499, n500, n501, n502, n503, n504, n505;
  wire n506, n507, n508, n509, n510, n511, n512, n513;
  wire n514, n515, n516, n517, n518, n519, n520, n521;
  wire n522, n523, n524, n525, n526, n527, n528, n529;
  wire n530, n531, n532, n533, n534, n535, n536, n537;
  wire n538, n539, n540, n541, n542, n543, n544, n545;
  wire n546, n547, n548, n549, n550, n551, n552, n553;
  wire n554, n555, n556, n557, n558, n559, n560, n561;
  wire n562, n563, n564, n565, n566, n567, n568, n569;
  wire n570, n571, n572, n573, n574, n575, n576, n577;
  wire n578, n579, n580, n581, n582, n583, n584, n585;
  wire n586, n587, n588, n589, n590, n591, n592, n593;
  wire n594, n595, n596, n597, n598, n599, n600, n601;
  wire n602, n603, n604, n605, n606, n607, n608, n609;
  wire n610, n611, n612, n613, n614, n615, n616, n617;
  wire n618, n619, n620, n621, n622, n623, n624, n625;
  wire n626, n627, n628, n629, n630, n631, n632, n633;
  wire n634, n635, n636, n637, n638, n639, n640, n641;
  wire n642, n643, n644, n645, n646, n647, n648, n649;
  wire n650, n651, n652, n653, n654, n655, n656, n657;
  wire n658, n659, n660, n661, n662, n663, n664, n665;
  wire n666, n667, n668, n669, n670, n671, n672, n673;
  wire n674, n675, n676, n677, n678, n679, n680, n681;
  wire n682, n683, n684, n685, n686, n687, n688, n689;
  wire n690, n691, n692, n693, n694, n695, n696, n697;
  wire n698, n699, n700, n701, n702, n703, n704, n705;
  wire n706, n707, n708, n709, n710, n711, n712, n713;
  wire n714, n715, n716, n717, n718, n719, n720, n721;
  wire n722, n723, n725, n726, n727, n728, n729, n730;
  wire n731, n732, n733, n734, n735, n736, n737, n738;
  wire n739, n740, n741, n742, n743, n744, n745, n746;
  wire n747, n748, n749, n750, n751, n752, n753, n754;
  wire n755, n756, n757, n758, n759, n760, n761, n762;
  wire n763, n764, n765, n766, n767, n768, n769, n770;
  wire n771, n772, n773, n774, n775, n776, n777, n778;
  wire n779, n780, n781, n782, n783, n784, n785, n786;
  wire n787, n788, n789, n790, n791, n792, n793, n794;
  wire n795, n796, n797, n798, n799, n800, n801, n802;
  wire n803, n804, n805, n806, n807, n808, n809, n810;
  wire n811, n812, n813, n814, n815, n816, n817, n818;
  wire n819, n820, n821, n822, n823, n824, n825, n826;
  wire n827, n828, n829, n830, n831, n832, n833, n834;
  wire n835, n836, n837, n838, n839, n840, n841, n842;
  wire n843, n844, n845, n846, n847, n848, n849, n850;
  wire n851, n852, n853, n854, n855, n856, n857, n858;
  wire n859, n860, n861, n862, n863, n864, n865, n866;
  wire n867, n868, n869, n870, n871, n872, n873, n874;
  wire n875, n876, n877, n878, n879, n880, n881, n882;
  wire n883, n884, n885, n886, n887, n888, n889, n890;
  wire n891, n892, n893, n894, n895, n896, n897, n898;
  wire n899, n900, n901, n902, n903, n904, n905, n906;
  wire n907, n908, n909, n910, n911, n912, n913, n914;
  wire n915, n916, n917, n918, n919, n920, n921, n922;
  wire n923, n924, n925, n926, n927, n928, n929, n930;
  wire n931, n932, n933, n934, n935, n936, n937, n938;
  wire n939, n940, n941, n942, n943, n944, n945, n946;
  wire n947, n948, n949, n950, n951, n952, n953, n954;
  wire n955, n956, n957, n958, n959, n960, n961, n962;
  wire n963, n964, n965, n966, n967, n968, n969, n970;
  wire n971, n972, n973, n974, n975, n976, n977, n978;
  wire n979, n980, n981, n982, n983, n984, n985, n986;
  wire n987, n988, n989, n990, n991, n992, n993, n994;
  wire n995, n996, n997, n998, n999, n1000, n1001, n1002;
  wire n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010;
  wire n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  wire n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  wire n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  wire n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  wire n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050;
  wire n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058;
  wire n1059, n1060, n1061, n1062, n1064, n1065, n1066, n1067;
  wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
  wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
  wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
  wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
  wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
  wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
  wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
  wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
  wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
  wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
  wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
  wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
  wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
  wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
  wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
  wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
  wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
  wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
  wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
  wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
  wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
  wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
  wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
  wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
  wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
  wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
  wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
  wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
  wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
  wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
  wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
  wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
  wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
  wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
  wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
  wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
  wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
  wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
  wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
  wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
  wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
  wire n1396, n1397, n1398, n1399, n1401, n1402, n1403, n1404;
  wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
  wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
  wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
  wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
  wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
  wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
  wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
  wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
  wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
  wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
  wire n1485, n1486, n1487, n1488, n1489, n1491, n1492, n1493;
  wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
  wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
  wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
  wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
  wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
  wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
  wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
  wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
  wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
  wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
  wire n1574, n1575, n1576, n1577, n1578, n1579, n1581, n1582;
  wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
  wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
  wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
  wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
  wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
  wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
  wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
  wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
  wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
  wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
  wire n1663, n1664, n1665, n1666, n1668, n1669, n1670, n1671;
  wire n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679;
  wire n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687;
  wire n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695;
  wire n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703;
  wire n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711;
  wire n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719;
  wire n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727;
  wire n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735;
  wire n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743;
  wire n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751;
  wire n1752, n1753, n1755, n1756, n1757, n1758, n1759, n1760;
  wire n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768;
  wire n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776;
  wire n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784;
  wire n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792;
  wire n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800;
  wire n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808;
  wire n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816;
  wire n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824;
  wire n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832;
  wire n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840;
  wire n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849;
  wire n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857;
  wire n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865;
  wire n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873;
  wire n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881;
  wire n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889;
  wire n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897;
  wire n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905;
  wire n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913;
  wire n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921;
  wire n1922, n1923, n1924, n1925, n1926, n1928, n1929, n1930;
  wire n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938;
  wire n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946;
  wire n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954;
  wire n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;
  wire n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970;
  wire n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978;
  wire n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986;
  wire n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994;
  wire n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002;
  wire n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010;
  wire n2011, n2012, n2014, n2015, n2016, n2017, n2018, n2019;
  wire n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027;
  wire n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035;
  wire n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043;
  wire n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051;
  wire n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059;
  wire n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067;
  wire n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075;
  wire n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083;
  wire n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091;
  wire n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2100;
  wire n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108;
  wire n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116;
  wire n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124;
  wire n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132;
  wire n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140;
  wire n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
  wire n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156;
  wire n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164;
  wire n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172;
  wire n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180;
  wire n2181, n2182, n2183, n2184, n2186, n2187, n2188, n2189;
  wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197;
  wire n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
  wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
  wire n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
  wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
  wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237;
  wire n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245;
  wire n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253;
  wire n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
  wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
  wire n2270, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
  wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
  wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
  wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
  wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
  wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
  wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
  wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
  wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
  wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
  wire n2351, n2352, n2353, n2354, n2355, n2356, n2358, n2359;
  wire n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367;
  wire n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375;
  wire n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383;
  wire n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391;
  wire n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399;
  wire n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407;
  wire n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415;
  wire n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423;
  wire n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431;
  wire n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439;
  wire n2440, n2441, n2442, n2444, n2445, n2446, n2447, n2448;
  wire n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456;
  wire n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464;
  wire n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472;
  wire n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480;
  wire n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488;
  wire n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496;
  wire n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504;
  wire n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512;
  wire n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520;
  wire n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528;
  wire n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537;
  wire n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545;
  wire n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553;
  wire n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561;
  wire n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569;
  wire n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577;
  wire n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585;
  wire n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593;
  wire n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601;
  wire n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609;
  wire n2610, n2611, n2612, n2613, n2614, n2616, n2617, n2618;
  wire n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626;
  wire n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634;
  wire n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642;
  wire n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650;
  wire n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658;
  wire n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666;
  wire n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674;
  wire n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682;
  wire n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690;
  wire n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698;
  wire n2699, n2700, n2702, n2703, n2704, n2705, n2706, n2707;
  wire n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715;
  wire n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723;
  wire n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731;
  wire n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739;
  wire n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747;
  wire n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755;
  wire n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763;
  wire n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771;
  wire n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779;
  wire n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2788;
  wire n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796;
  wire n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804;
  wire n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812;
  wire n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820;
  wire n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828;
  wire n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836;
  wire n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844;
  wire n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852;
  wire n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860;
  wire n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868;
  wire n2869, n2870, n2871, n2872, n2874, n2875, n2876, n2877;
  wire n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885;
  wire n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893;
  wire n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901;
  wire n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909;
  wire n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917;
  wire n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925;
  wire n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933;
  wire n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941;
  wire n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949;
  wire n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957;
  wire n2958, n2960, n2961, n2962, n2963, n2964, n2965, n2966;
  wire n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974;
  wire n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982;
  wire n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990;
  wire n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998;
  wire n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006;
  wire n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014;
  wire n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022;
  wire n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030;
  wire n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038;
  wire n3039, n3040, n3041, n3042, n3043, n3044, n3046, n3047;
  wire n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055;
  wire n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063;
  wire n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071;
  wire n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079;
  wire n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087;
  wire n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095;
  wire n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103;
  wire n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111;
  wire n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119;
  wire n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127;
  wire n3128, n3129, n3130, n3132, n3133, n3134, n3135, n3136;
  wire n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144;
  wire n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152;
  wire n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160;
  wire n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168;
  wire n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176;
  wire n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184;
  wire n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192;
  wire n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200;
  wire n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208;
  wire n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216;
  wire n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225;
  wire n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233;
  wire n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241;
  wire n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249;
  wire n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257;
  wire n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265;
  wire n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273;
  wire n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281;
  wire n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289;
  wire n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297;
  wire n3298, n3299, n3300, n3301, n3302, n3304, n3305, n3306;
  wire n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314;
  wire n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322;
  wire n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330;
  wire n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338;
  wire n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346;
  wire n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354;
  wire n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362;
  wire n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370;
  wire n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378;
  wire n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386;
  wire n3387, n3388, n3390, n3391, n3392, n3393, n3394, n3395;
  wire n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403;
  wire n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411;
  wire n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419;
  wire n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427;
  wire n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435;
  wire n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443;
  wire n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451;
  wire n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459;
  wire n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467;
  wire n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3476;
  wire n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484;
  wire n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492;
  wire n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500;
  wire n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508;
  wire n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516;
  wire n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524;
  wire n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532;
  wire n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540;
  wire n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548;
  wire n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556;
  wire n3557, n3558, n3559, n3560, n3562, n3563, n3564, n3565;
  wire n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573;
  wire n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581;
  wire n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589;
  wire n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597;
  wire n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605;
  wire n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613;
  wire n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621;
  wire n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629;
  wire n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637;
  wire n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645;
  wire n3646, n3648, n3649, n3650, n3651, n3652, n3653, n3654;
  wire n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662;
  wire n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670;
  wire n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678;
  wire n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686;
  wire n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694;
  wire n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702;
  wire n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710;
  wire n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718;
  wire n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726;
  wire n3727, n3728, n3729, n3730, n3731, n3732, n3734, n3735;
  wire n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743;
  wire n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751;
  wire n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759;
  wire n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767;
  wire n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775;
  wire n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783;
  wire n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791;
  wire n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799;
  wire n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807;
  wire n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815;
  wire n3816, n3817, n3818, n3820, n3821, n3822, n3823, n3824;
  wire n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832;
  wire n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840;
  wire n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848;
  wire n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856;
  wire n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864;
  wire n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872;
  wire n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880;
  wire n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888;
  wire n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896;
  wire n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904;
  wire n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913;
  wire n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921;
  wire n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929;
  wire n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937;
  wire n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945;
  wire n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953;
  wire n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961;
  wire n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969;
  wire n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977;
  wire n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985;
  wire n3986, n3987, n3988, n3989, n3990, n3992, n3993, n3994;
  wire n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002;
  wire n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010;
  wire n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018;
  wire n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026;
  wire n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034;
  wire n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042;
  wire n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050;
  wire n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058;
  wire n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066;
  wire n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074;
  wire n4075, n4076, n4078, n4079, n4080, n4081, n4082, n4083;
  wire n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091;
  wire n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099;
  wire n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107;
  wire n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115;
  wire n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123;
  wire n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131;
  wire n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139;
  wire n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147;
  wire n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155;
  wire n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4164;
  wire n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172;
  wire n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180;
  wire n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188;
  wire n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196;
  wire n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204;
  wire n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212;
  wire n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220;
  wire n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228;
  wire n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236;
  wire n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244;
  wire n4245, n4246, n4247, n4248, n4250, n4251, n4252, n4253;
  wire n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261;
  wire n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269;
  wire n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277;
  wire n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285;
  wire n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293;
  wire n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301;
  wire n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309;
  wire n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317;
  wire n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325;
  wire n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333;
  wire n4334, n4336, n4337, n4338, n4339, n4340, n4341, n4342;
  wire n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350;
  wire n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358;
  wire n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366;
  wire n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374;
  wire n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382;
  wire n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390;
  wire n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398;
  wire n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406;
  wire n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414;
  wire n4415, n4416, n4417, n4418, n4419, n4420, n4422, n4423;
  wire n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431;
  wire n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439;
  wire n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447;
  wire n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455;
  wire n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463;
  wire n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471;
  wire n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479;
  wire n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487;
  wire n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495;
  wire n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503;
  wire n4504, n4505, n4506, n4508, n4509, n4510, n4511, n4512;
  wire n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520;
  wire n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528;
  wire n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536;
  wire n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544;
  wire n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552;
  wire n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560;
  wire n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568;
  wire n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576;
  wire n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584;
  wire n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592;
  wire n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601;
  wire n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609;
  wire n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617;
  wire n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625;
  wire n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633;
  wire n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641;
  wire n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649;
  wire n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657;
  wire n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665;
  wire n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673;
  wire n4674, n4675, n4676, n4677, n4678, n4680, n4681, n4682;
  wire n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690;
  wire n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698;
  wire n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706;
  wire n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714;
  wire n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722;
  wire n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730;
  wire n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738;
  wire n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746;
  wire n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754;
  wire n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762;
  wire n4763, n4764, n4766, n4767, n4768, n4769, n4770, n4771;
  wire n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779;
  wire n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787;
  wire n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795;
  wire n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803;
  wire n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811;
  wire n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819;
  wire n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827;
  wire n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835;
  wire n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843;
  wire n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4852;
  wire n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860;
  wire n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868;
  wire n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876;
  wire n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884;
  wire n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892;
  wire n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900;
  wire n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908;
  wire n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916;
  wire n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924;
  wire n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932;
  wire n4933, n4934, n4935, n4936, n4938, n4939, n4940, n4941;
  wire n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949;
  wire n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957;
  wire n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965;
  wire n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973;
  wire n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981;
  wire n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989;
  wire n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997;
  wire n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005;
  wire n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013;
  wire n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021;
  wire n5022, n5024, n5025, n5026, n5027, n5028, n5029, n5030;
  wire n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038;
  wire n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046;
  wire n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054;
  wire n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062;
  wire n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070;
  wire n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078;
  wire n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086;
  wire n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094;
  wire n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102;
  wire n5103, n5104, n5105, n5106, n5107, n5108, n5110, n5111;
  wire n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119;
  wire n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127;
  wire n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135;
  wire n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143;
  wire n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151;
  wire n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159;
  wire n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167;
  wire n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175;
  wire n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183;
  wire n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191;
  wire n5192, n5193, n5194, n5196, n5197, n5198, n5199, n5200;
  wire n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208;
  wire n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216;
  wire n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224;
  wire n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232;
  wire n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240;
  wire n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248;
  wire n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256;
  wire n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264;
  wire n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272;
  wire n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280;
  wire n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289;
  wire n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297;
  wire n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305;
  wire n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313;
  wire n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321;
  wire n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329;
  wire n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337;
  wire n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345;
  wire n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353;
  wire n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361;
  wire n5362, n5363, n5364, n5365, n5366, n5368, n5369, n5370;
  wire n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378;
  wire n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386;
  wire n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394;
  wire n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402;
  wire n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410;
  wire n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418;
  wire n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426;
  wire n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434;
  wire n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442;
  wire n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450;
  wire n5451, n5452, n5454, n5455, n5456, n5457, n5458, n5459;
  wire n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467;
  wire n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475;
  wire n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483;
  wire n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491;
  wire n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499;
  wire n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507;
  wire n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515;
  wire n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523;
  wire n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531;
  wire n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5540;
  wire n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548;
  wire n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556;
  wire n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564;
  wire n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572;
  wire n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580;
  wire n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588;
  wire n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596;
  wire n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604;
  wire n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612;
  wire n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620;
  wire n5621, n5622, n5623, n5624, n5626, n5627, n5628, n5629;
  wire n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637;
  wire n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645;
  wire n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653;
  wire n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661;
  wire n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669;
  wire n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677;
  wire n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685;
  wire n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693;
  wire n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701;
  wire n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709;
  wire n5710, n5712, n5713, n5714, n5715, n5716, n5717, n5718;
  wire n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726;
  wire n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734;
  wire n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742;
  wire n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750;
  wire n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758;
  wire n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766;
  wire n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774;
  wire n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782;
  wire n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790;
  wire n5791, n5792, n5793, n5794, n5795, n5796, n5798, n5799;
  wire n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807;
  wire n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815;
  wire n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823;
  wire n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831;
  wire n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839;
  wire n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847;
  wire n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855;
  wire n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863;
  wire n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871;
  wire n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879;
  wire n5880, n5881, n5882, n5884, n5885, n5886, n5887, n5888;
  wire n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896;
  wire n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904;
  wire n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912;
  wire n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920;
  wire n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928;
  wire n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936;
  wire n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944;
  wire n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952;
  wire n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960;
  wire n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968;
  wire n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977;
  wire n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985;
  wire n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993;
  wire n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001;
  wire n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009;
  wire n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017;
  wire n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025;
  wire n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033;
  wire n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041;
  wire n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049;
  wire n6050, n6051, n6052, n6053, n6054, n6056, n6057, n6058;
  wire n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066;
  wire n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074;
  wire n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082;
  wire n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090;
  wire n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098;
  wire n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106;
  wire n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114;
  wire n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122;
  wire n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130;
  wire n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138;
  wire n6139, n6140, n6142, n6143, n6144, n6145, n6146, n6147;
  wire n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155;
  wire n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163;
  wire n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171;
  wire n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179;
  wire n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187;
  wire n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195;
  wire n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203;
  wire n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211;
  wire n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219;
  wire n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6228;
  wire n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236;
  wire n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244;
  wire n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252;
  wire n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260;
  wire n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268;
  wire n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276;
  wire n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284;
  wire n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292;
  wire n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300;
  wire n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308;
  wire n6309, n6310, n6311, n6312, n6314, n6315, n6316, n6317;
  wire n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325;
  wire n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333;
  wire n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341;
  wire n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349;
  wire n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357;
  wire n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365;
  wire n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373;
  wire n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381;
  wire n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389;
  wire n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397;
  wire n6398, n6400, n6401, n6402, n6403, n6404, n6405, n6406;
  wire n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414;
  wire n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422;
  wire n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430;
  wire n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438;
  wire n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446;
  wire n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454;
  wire n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462;
  wire n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470;
  wire n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478;
  wire n6479, n6480, n6481, n6482, n6483, n6484, n6486, n6487;
  wire n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495;
  wire n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503;
  wire n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511;
  wire n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519;
  wire n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527;
  wire n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535;
  wire n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543;
  wire n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551;
  wire n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559;
  wire n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567;
  wire n6568, n6569, n6570, n6572, n6573, n6574, n6575, n6576;
  wire n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584;
  wire n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592;
  wire n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600;
  wire n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608;
  wire n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616;
  wire n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624;
  wire n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632;
  wire n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640;
  wire n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648;
  wire n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656;
  wire n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665;
  wire n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673;
  wire n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681;
  wire n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689;
  wire n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697;
  wire n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705;
  wire n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713;
  wire n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721;
  wire n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729;
  wire n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737;
  wire n6738, n6739, n6740, n6741, n6742, n6744, n6745, n6746;
  wire n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754;
  wire n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762;
  wire n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770;
  wire n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778;
  wire n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786;
  wire n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794;
  wire n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802;
  wire n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810;
  wire n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818;
  wire n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826;
  wire n6827, n6828, n6830, n6831, n6832, n6833, n6834, n6835;
  wire n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843;
  wire n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851;
  wire n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859;
  wire n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867;
  wire n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875;
  wire n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883;
  wire n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891;
  wire n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899;
  wire n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907;
  wire n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6916;
  wire n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924;
  wire n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932;
  wire n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940;
  wire n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948;
  wire n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956;
  wire n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964;
  wire n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972;
  wire n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980;
  wire n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988;
  wire n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996;
  wire n6997, n6998, n6999, n7000, n7002, n7003, n7004, n7005;
  wire n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013;
  wire n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021;
  wire n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029;
  wire n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037;
  wire n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045;
  wire n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053;
  wire n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061;
  wire n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069;
  wire n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077;
  wire n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085;
  wire n7086, n7088, n7089, n7090, n7091, n7092, n7093, n7094;
  wire n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102;
  wire n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110;
  wire n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118;
  wire n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126;
  wire n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134;
  wire n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142;
  wire n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150;
  wire n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158;
  wire n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166;
  wire n7167, n7168, n7169, n7170, n7171, n7172, n7174, n7175;
  wire n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183;
  wire n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191;
  wire n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199;
  wire n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207;
  wire n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215;
  wire n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223;
  wire n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231;
  wire n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239;
  wire n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247;
  wire n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255;
  wire n7256, n7257, n7258, n7260, n7261, n7262, n7263, n7264;
  wire n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272;
  wire n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280;
  wire n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288;
  wire n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296;
  wire n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304;
  wire n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312;
  wire n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320;
  wire n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328;
  wire n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336;
  wire n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344;
  wire n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353;
  wire n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361;
  wire n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369;
  wire n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377;
  wire n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385;
  wire n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393;
  wire n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401;
  wire n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409;
  wire n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417;
  wire n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425;
  wire n7426, n7427, n7428, n7429, n7430, n7432, n7433, n7434;
  wire n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442;
  wire n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450;
  wire n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458;
  wire n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466;
  wire n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474;
  wire n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482;
  wire n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490;
  wire n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498;
  wire n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506;
  wire n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514;
  wire n7515, n7516, n7518, n7519, n7520, n7521, n7522, n7523;
  wire n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531;
  wire n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539;
  wire n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547;
  wire n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555;
  wire n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563;
  wire n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571;
  wire n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579;
  wire n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587;
  wire n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595;
  wire n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7604;
  wire n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612;
  wire n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620;
  wire n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628;
  wire n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636;
  wire n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644;
  wire n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652;
  wire n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660;
  wire n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668;
  wire n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676;
  wire n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684;
  wire n7685, n7686, n7687, n7688, n7690, n7691, n7692, n7693;
  wire n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701;
  wire n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709;
  wire n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717;
  wire n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725;
  wire n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733;
  wire n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741;
  wire n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749;
  wire n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757;
  wire n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765;
  wire n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773;
  wire n7774, n7776, n7777, n7778, n7779, n7780, n7781, n7782;
  wire n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790;
  wire n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798;
  wire n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806;
  wire n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814;
  wire n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822;
  wire n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830;
  wire n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838;
  wire n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846;
  wire n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854;
  wire n7855, n7856, n7857, n7858, n7859, n7860, n7862, n7863;
  wire n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871;
  wire n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879;
  wire n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887;
  wire n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895;
  wire n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903;
  wire n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911;
  wire n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919;
  wire n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927;
  wire n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935;
  wire n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943;
  wire n7944, n7945, n7946, n7948, n7949, n7950, n7951, n7952;
  wire n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960;
  wire n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968;
  wire n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976;
  wire n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984;
  wire n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992;
  wire n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000;
  wire n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008;
  wire n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016;
  wire n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024;
  wire n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032;
  wire n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041;
  wire n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049;
  wire n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057;
  wire n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065;
  wire n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073;
  wire n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081;
  wire n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089;
  wire n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097;
  wire n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105;
  wire n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113;
  wire n8114, n8115, n8116, n8117, n8118, n8120, n8121, n8122;
  wire n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130;
  wire n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138;
  wire n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146;
  wire n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154;
  wire n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162;
  wire n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170;
  wire n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178;
  wire n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186;
  wire n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194;
  wire n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202;
  wire n8203, n8204, n8206, n8207, n8208, n8209, n8210, n8211;
  wire n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219;
  wire n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227;
  wire n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235;
  wire n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243;
  wire n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251;
  wire n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259;
  wire n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267;
  wire n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275;
  wire n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283;
  wire n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8292;
  wire n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300;
  wire n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308;
  wire n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316;
  wire n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324;
  wire n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332;
  wire n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340;
  wire n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348;
  wire n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356;
  wire n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364;
  wire n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372;
  wire n8373, n8374, n8375, n8376, n8378, n8379, n8380, n8381;
  wire n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389;
  wire n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397;
  wire n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405;
  wire n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413;
  wire n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421;
  wire n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429;
  wire n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437;
  wire n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445;
  wire n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453;
  wire n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461;
  wire n8462, n8464, n8465, n8466, n8467, n8468, n8469, n8470;
  wire n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478;
  wire n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486;
  wire n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494;
  wire n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502;
  wire n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510;
  wire n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518;
  wire n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526;
  wire n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534;
  wire n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542;
  wire n8543, n8544, n8545, n8546, n8547, n8548, n8550, n8551;
  wire n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559;
  wire n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567;
  wire n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575;
  wire n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583;
  wire n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591;
  wire n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599;
  wire n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607;
  wire n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615;
  wire n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623;
  wire n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631;
  wire n8632, n8633, n8634, n8636, n8637, n8638, n8639, n8640;
  wire n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648;
  wire n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656;
  wire n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664;
  wire n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672;
  wire n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680;
  wire n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688;
  wire n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696;
  wire n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704;
  wire n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712;
  wire n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720;
  wire n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729;
  wire n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737;
  wire n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745;
  wire n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753;
  wire n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761;
  wire n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769;
  wire n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777;
  wire n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785;
  wire n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793;
  wire n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801;
  wire n8802, n8803, n8804, n8805, n8806, n8808, n8809, n8810;
  wire n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818;
  wire n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826;
  wire n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834;
  wire n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842;
  wire n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850;
  wire n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858;
  wire n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866;
  wire n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874;
  wire n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882;
  wire n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890;
  wire n8891, n8892, n8894, n8895, n8896, n8897, n8898, n8899;
  wire n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907;
  wire n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915;
  wire n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923;
  wire n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931;
  wire n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939;
  wire n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947;
  wire n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955;
  wire n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963;
  wire n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971;
  wire n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8980;
  wire n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988;
  wire n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996;
  wire n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004;
  wire n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012;
  wire n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020;
  wire n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028;
  wire n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036;
  wire n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044;
  wire n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052;
  wire n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060;
  wire n9061, n9062, n9063, n9064, n9066, n9067, n9068, n9069;
  wire n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077;
  wire n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085;
  wire n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093;
  wire n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101;
  wire n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109;
  wire n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117;
  wire n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125;
  wire n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133;
  wire n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141;
  wire n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149;
  wire n9150, n9152, n9153, n9154, n9155, n9156, n9157, n9158;
  wire n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166;
  wire n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174;
  wire n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182;
  wire n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190;
  wire n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198;
  wire n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206;
  wire n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214;
  wire n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222;
  wire n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230;
  wire n9231, n9232, n9233, n9234, n9235, n9236, n9238, n9239;
  wire n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247;
  wire n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255;
  wire n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263;
  wire n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271;
  wire n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279;
  wire n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287;
  wire n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295;
  wire n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303;
  wire n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311;
  wire n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319;
  wire n9320, n9321, n9322, n9324, n9325, n9326, n9327, n9328;
  wire n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336;
  wire n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344;
  wire n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352;
  wire n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360;
  wire n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368;
  wire n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376;
  wire n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384;
  wire n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392;
  wire n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400;
  wire n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408;
  wire n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417;
  wire n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425;
  wire n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433;
  wire n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441;
  wire n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449;
  wire n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457;
  wire n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465;
  wire n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473;
  wire n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481;
  wire n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489;
  wire n9490, n9491, n9492, n9493, n9494, n9496, n9497, n9498;
  wire n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506;
  wire n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514;
  wire n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522;
  wire n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530;
  wire n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538;
  wire n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546;
  wire n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554;
  wire n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562;
  wire n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570;
  wire n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578;
  wire n9579, n9580, n9582, n9583, n9584, n9585, n9586, n9587;
  wire n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595;
  wire n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603;
  wire n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611;
  wire n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619;
  wire n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627;
  wire n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635;
  wire n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643;
  wire n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651;
  wire n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659;
  wire n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9668;
  wire n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676;
  wire n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684;
  wire n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692;
  wire n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700;
  wire n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708;
  wire n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716;
  wire n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724;
  wire n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732;
  wire n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740;
  wire n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748;
  wire n9749, n9750, n9751, n9752, n9754, n9755, n9756, n9757;
  wire n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765;
  wire n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773;
  wire n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781;
  wire n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789;
  wire n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797;
  wire n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805;
  wire n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813;
  wire n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821;
  wire n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829;
  wire n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837;
  wire n9838, n9840, n9841, n9842, n9843, n9844, n9845, n9846;
  wire n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854;
  wire n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862;
  wire n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870;
  wire n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878;
  wire n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886;
  wire n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894;
  wire n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902;
  wire n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910;
  wire n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918;
  wire n9919, n9920, n9921, n9922, n9923, n9924, n9926, n9927;
  wire n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935;
  wire n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943;
  wire n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951;
  wire n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959;
  wire n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967;
  wire n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975;
  wire n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983;
  wire n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991;
  wire n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999;
  wire n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007;
  wire n10008, n10009, n10010, n10012, n10013, n10014, n10015, n10016;
  wire n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024;
  wire n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032;
  wire n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040;
  wire n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048;
  wire n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056;
  wire n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064;
  wire n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072;
  wire n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080;
  wire n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088;
  wire n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096;
  wire n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105;
  wire n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113;
  wire n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121;
  wire n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129;
  wire n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137;
  wire n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145;
  wire n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153;
  wire n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161;
  wire n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169;
  wire n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177;
  wire n10178, n10179, n10180, n10181, n10182, n10184, n10185, n10186;
  wire n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194;
  wire n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202;
  wire n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210;
  wire n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218;
  wire n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226;
  wire n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234;
  wire n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242;
  wire n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250;
  wire n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258;
  wire n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266;
  wire n10267, n10268, n10270, n10271, n10272, n10273, n10274, n10275;
  wire n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283;
  wire n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291;
  wire n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299;
  wire n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307;
  wire n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315;
  wire n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323;
  wire n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331;
  wire n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339;
  wire n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347;
  wire n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10356;
  wire n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364;
  wire n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372;
  wire n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380;
  wire n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388;
  wire n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396;
  wire n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404;
  wire n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412;
  wire n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420;
  wire n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428;
  wire n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436;
  wire n10437, n10438, n10439, n10440, n10442, n10443, n10444, n10445;
  wire n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453;
  wire n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461;
  wire n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469;
  wire n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477;
  wire n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485;
  wire n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493;
  wire n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501;
  wire n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509;
  wire n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517;
  wire n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525;
  wire n10526, n10528, n10529, n10530, n10531, n10532, n10533, n10534;
  wire n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542;
  wire n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550;
  wire n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558;
  wire n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566;
  wire n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574;
  wire n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582;
  wire n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590;
  wire n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598;
  wire n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606;
  wire n10607, n10608, n10609, n10610, n10611, n10612, n10614, n10615;
  wire n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623;
  wire n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631;
  wire n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639;
  wire n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647;
  wire n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655;
  wire n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663;
  wire n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671;
  wire n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679;
  wire n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687;
  wire n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695;
  wire n10696, n10697, n10698, n10700, n10701, n10702, n10703, n10704;
  wire n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712;
  wire n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720;
  wire n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728;
  wire n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736;
  wire n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744;
  wire n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752;
  wire n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760;
  wire n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768;
  wire n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776;
  wire n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784;
  wire n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793;
  wire n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801;
  wire n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809;
  wire n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817;
  wire n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825;
  wire n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833;
  wire n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841;
  wire n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849;
  wire n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857;
  wire n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865;
  wire n10866, n10867, n10868, n10869, n10870, n10872, n10873, n10874;
  wire n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882;
  wire n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890;
  wire n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898;
  wire n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906;
  wire n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914;
  wire n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922;
  wire n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930;
  wire n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938;
  wire n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946;
  wire n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954;
  wire n10955, n10956, n10958, n10959, n10960, n10961, n10962, n10963;
  wire n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971;
  wire n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979;
  wire n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987;
  wire n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995;
  wire n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003;
  wire n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011;
  wire n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019;
  wire n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027;
  wire n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035;
  wire n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11044;
  wire n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052;
  wire n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060;
  wire n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068;
  wire n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076;
  wire n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084;
  wire n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092;
  wire n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100;
  wire n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108;
  wire n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116;
  wire n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124;
  wire n11125, n11126, n11127, n11128, n11130, n11131, n11132, n11133;
  wire n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141;
  wire n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149;
  wire n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157;
  wire n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165;
  wire n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173;
  wire n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181;
  wire n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189;
  wire n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197;
  wire n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205;
  wire n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213;
  wire n11214, n11216, n11217, n11218, n11219, n11220, n11221, n11222;
  wire n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230;
  wire n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238;
  wire n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246;
  wire n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254;
  wire n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262;
  wire n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270;
  wire n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278;
  wire n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286;
  wire n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294;
  wire n11295, n11296, n11297, n11298, n11299, n11300, n11302, n11303;
  wire n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311;
  wire n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319;
  wire n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327;
  wire n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335;
  wire n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343;
  wire n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351;
  wire n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359;
  wire n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367;
  wire n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375;
  wire n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383;
  wire n11384, n11385, n11386, n11388, n11389, n11390, n11391, n11392;
  wire n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400;
  wire n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408;
  wire n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416;
  wire n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424;
  wire n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432;
  wire n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440;
  wire n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448;
  wire n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456;
  wire n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464;
  wire n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472;
  wire n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481;
  wire n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489;
  wire n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497;
  wire n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505;
  wire n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513;
  wire n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521;
  wire n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529;
  wire n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537;
  wire n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545;
  wire n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553;
  wire n11554, n11555, n11556, n11557, n11558, n11560, n11561, n11562;
  wire n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570;
  wire n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578;
  wire n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586;
  wire n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594;
  wire n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602;
  wire n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610;
  wire n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618;
  wire n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626;
  wire n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634;
  wire n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642;
  wire n11643, n11644, n11646, n11647, n11648, n11649, n11650, n11651;
  wire n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659;
  wire n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667;
  wire n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675;
  wire n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683;
  wire n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691;
  wire n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699;
  wire n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707;
  wire n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715;
  wire n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723;
  wire n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11732;
  wire n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740;
  wire n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748;
  wire n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756;
  wire n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764;
  wire n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772;
  wire n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780;
  wire n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788;
  wire n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796;
  wire n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804;
  wire n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812;
  wire n11813, n11814, n11815, n11816, n11818, n11819, n11820, n11821;
  wire n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829;
  wire n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837;
  wire n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845;
  wire n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853;
  wire n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861;
  wire n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869;
  wire n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877;
  wire n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885;
  wire n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893;
  wire n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901;
  wire n11902, n11904, n11905, n11906, n11907, n11908, n11909, n11910;
  wire n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918;
  wire n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926;
  wire n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934;
  wire n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942;
  wire n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950;
  wire n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958;
  wire n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966;
  wire n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974;
  wire n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982;
  wire n11983, n11984, n11985, n11986, n11987, n11988, n11990, n11991;
  wire n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999;
  wire n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007;
  wire n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015;
  wire n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023;
  wire n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031;
  wire n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039;
  wire n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047;
  wire n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055;
  wire n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063;
  wire n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071;
  wire n12072, n12073, n12074, n12076, n12077, n12078, n12079, n12080;
  wire n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088;
  wire n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096;
  wire n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104;
  wire n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112;
  wire n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120;
  wire n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128;
  wire n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136;
  wire n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144;
  wire n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152;
  wire n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160;
  wire n_3, n_5, n_6, n_9, n_10, n_11, n_14, n_15;
  wire n_17, n_18, n_22, n_23, n_24, n_25, n_28, n_29;
  wire n_31, n_32, n_36, n_37, n_38, n_39, n_42, n_43;
  wire n_45, n_46, n_50, n_51, n_52, n_53, n_56, n_57;
  wire n_59, n_60, n_64, n_65, n_66, n_67, n_70, n_71;
  wire n_73, n_74, n_78, n_79, n_80, n_81, n_84, n_85;
  wire n_87, n_88, n_92, n_93, n_94, n_95, n_98, n_99;
  wire n_101, n_102, n_106, n_107, n_108, n_109, n_112, n_113;
  wire n_115, n_116, n_120, n_121, n_122, n_123, n_126, n_127;
  wire n_129, n_130, n_134, n_135, n_136, n_137, n_140, n_141;
  wire n_143, n_144, n_148, n_149, n_150, n_151, n_154, n_155;
  wire n_157, n_158, n_162, n_163, n_164, n_165, n_168, n_169;
  wire n_171, n_172, n_176, n_177, n_178, n_179, n_182, n_183;
  wire n_185, n_186, n_190, n_191, n_192, n_193, n_196, n_197;
  wire n_199, n_200, n_204, n_205, n_206, n_207, n_210, n_211;
  wire n_213, n_214, n_218, n_219, n_220, n_221, n_224, n_225;
  wire n_227, n_228, n_232, n_233, n_234, n_235, n_238, n_239;
  wire n_241, n_242, n_246, n_247, n_248, n_249, n_252, n_253;
  wire n_255, n_256, n_260, n_261, n_262, n_263, n_266, n_267;
  wire n_269, n_270, n_274, n_275, n_276, n_277, n_280, n_281;
  wire n_283, n_284, n_288, n_289, n_290, n_291, n_294, n_295;
  wire n_297, n_298, n_302, n_303, n_304, n_305, n_308, n_309;
  wire n_311, n_312, n_316, n_317, n_318, n_319, n_322, n_323;
  wire n_325, n_326, n_330, n_331, n_332, n_333, n_336, n_337;
  wire n_339, n_340, n_344, n_345, n_346, n_347, n_350, n_351;
  wire n_353, n_354, n_358, n_359, n_360, n_361, n_364, n_365;
  wire n_367, n_368, n_372, n_373, n_374, n_375, n_378, n_379;
  wire n_381, n_382, n_386, n_387, n_388, n_389, n_392, n_393;
  wire n_395, n_396, n_400, n_401, n_402, n_403, n_406, n_407;
  wire n_409, n_410, n_414, n_415, n_416, n_417, n_420, n_421;
  wire n_423, n_424, n_428, n_429, n_430, n_431, n_434, n_435;
  wire n_437, n_438, n_442, n_443, n_444, n_445, n_448, n_449;
  wire n_451, n_452, n_456, n_457, n_458, n_459, n_462, n_463;
  wire n_465, n_466, n_470, n_471, n_472, n_473, n_476, n_477;
  wire n_479, n_480, n_484, n_485, n_486, n_487, n_490, n_491;
  wire n_493, n_494, n_498, n_499, n_500, n_501, n_504, n_505;
  wire n_507, n_508, n_512, n_513, n_514, n_515, n_518, n_519;
  wire n_521, n_522, n_526, n_527, n_528, n_529, n_532, n_533;
  wire n_535, n_536, n_540, n_541, n_542, n_543, n_546, n_547;
  wire n_549, n_550, n_554, n_555, n_556, n_557, n_560, n_561;
  wire n_563, n_564, n_568, n_569, n_570, n_571, n_574, n_575;
  wire n_577, n_578, n_582, n_583, n_584, n_585, n_588, n_589;
  wire n_591, n_592, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672;
  wire n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704;
  wire n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784;
  wire n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792;
  wire n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800;
  wire n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808;
  wire n_809, n_810, n_811, n_812, n_813, n_814, n_815, n_816;
  wire n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840;
  wire n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848;
  wire n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864;
  wire n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872;
  wire n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880;
  wire n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896;
  wire n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904;
  wire n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936;
  wire n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944;
  wire n_945, n_946, n_947, n_948, n_949, n_950, n_951, n_952;
  wire n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960;
  wire n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968;
  wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
  wire n_977, n_978, n_979, n_980, n_981, n_982, n_983, n_984;
  wire n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016;
  wire n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048;
  wire n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088;
  wire n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096;
  wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104;
  wire n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112;
  wire n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120;
  wire n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128;
  wire n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152;
  wire n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184;
  wire n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272;
  wire n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280;
  wire n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288;
  wire n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320;
  wire n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336;
  wire n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344;
  wire n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
  wire n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360;
  wire n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368;
  wire n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376;
  wire n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408;
  wire n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416;
  wire n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424;
  wire n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432;
  wire n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440;
  wire n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448;
  wire n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456;
  wire n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464;
  wire n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472;
  wire n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480;
  wire n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488;
  wire n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496;
  wire n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504;
  wire n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512;
  wire n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520;
  wire n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528;
  wire n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536;
  wire n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544;
  wire n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552;
  wire n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568;
  wire n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576;
  wire n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600;
  wire n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608;
  wire n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616;
  wire n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624;
  wire n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632;
  wire n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648;
  wire n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656;
  wire n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664;
  wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672;
  wire n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680;
  wire n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728;
  wire n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736;
  wire n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744;
  wire n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752;
  wire n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
  wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872;
  wire n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880;
  wire n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888;
  wire n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896;
  wire n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920;
  wire n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928;
  wire n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936;
  wire n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984;
  wire n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992;
  wire n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016;
  wire n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040;
  wire n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048;
  wire n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056;
  wire n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064;
  wire n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072;
  wire n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080;
  wire n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088;
  wire n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096;
  wire n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104;
  wire n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112;
  wire n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120;
  wire n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128;
  wire n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136;
  wire n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144;
  wire n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152;
  wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
  wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
  wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176;
  wire n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184;
  wire n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192;
  wire n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200;
  wire n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224;
  wire n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232;
  wire n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240;
  wire n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248;
  wire n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256;
  wire n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264;
  wire n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272;
  wire n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280;
  wire n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288;
  wire n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296;
  wire n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304;
  wire n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312;
  wire n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320;
  wire n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328;
  wire n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336;
  wire n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344;
  wire n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352;
  wire n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360;
  wire n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368;
  wire n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376;
  wire n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384;
  wire n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392;
  wire n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400;
  wire n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408;
  wire n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416;
  wire n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424;
  wire n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432;
  wire n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440;
  wire n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448;
  wire n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456;
  wire n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464;
  wire n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472;
  wire n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480;
  wire n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488;
  wire n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496;
  wire n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504;
  wire n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512;
  wire n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520;
  wire n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528;
  wire n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536;
  wire n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544;
  wire n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552;
  wire n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560;
  wire n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568;
  wire n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576;
  wire n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584;
  wire n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592;
  wire n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600;
  wire n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608;
  wire n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616;
  wire n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624;
  wire n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632;
  wire n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640;
  wire n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648;
  wire n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656;
  wire n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664;
  wire n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
  wire n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680;
  wire n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688;
  wire n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696;
  wire n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704;
  wire n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712;
  wire n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744;
  wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
  wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
  wire n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768;
  wire n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776;
  wire n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784;
  wire n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792;
  wire n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800;
  wire n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808;
  wire n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816;
  wire n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824;
  wire n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832;
  wire n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840;
  wire n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848;
  wire n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856;
  wire n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864;
  wire n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872;
  wire n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880;
  wire n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888;
  wire n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896;
  wire n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904;
  wire n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912;
  wire n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920;
  wire n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928;
  wire n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936;
  wire n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944;
  wire n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952;
  wire n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960;
  wire n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968;
  wire n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976;
  wire n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984;
  wire n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992;
  wire n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000;
  wire n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008;
  wire n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016;
  wire n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024;
  wire n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032;
  wire n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040;
  wire n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048;
  wire n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056;
  wire n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064;
  wire n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072;
  wire n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080;
  wire n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088;
  wire n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096;
  wire n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104;
  wire n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112;
  wire n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120;
  wire n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128;
  wire n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136;
  wire n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144;
  wire n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152;
  wire n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160;
  wire n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168;
  wire n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176;
  wire n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184;
  wire n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192;
  wire n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200;
  wire n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208;
  wire n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216;
  wire n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224;
  wire n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232;
  wire n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240;
  wire n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248;
  wire n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256;
  wire n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264;
  wire n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272;
  wire n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280;
  wire n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288;
  wire n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296;
  wire n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304;
  wire n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312;
  wire n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320;
  wire n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328;
  wire n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336;
  wire n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344;
  wire n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352;
  wire n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360;
  wire n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368;
  wire n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376;
  wire n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384;
  wire n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392;
  wire n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400;
  wire n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408;
  wire n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416;
  wire n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424;
  wire n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432;
  wire n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440;
  wire n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448;
  wire n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456;
  wire n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464;
  wire n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472;
  wire n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480;
  wire n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488;
  wire n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496;
  wire n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504;
  wire n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512;
  wire n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520;
  wire n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528;
  wire n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536;
  wire n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544;
  wire n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552;
  wire n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560;
  wire n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568;
  wire n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576;
  wire n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584;
  wire n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592;
  wire n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600;
  wire n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608;
  wire n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616;
  wire n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624;
  wire n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632;
  wire n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640;
  wire n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648;
  wire n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656;
  wire n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664;
  wire n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672;
  wire n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680;
  wire n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688;
  wire n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696;
  wire n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704;
  wire n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712;
  wire n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720;
  wire n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728;
  wire n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736;
  wire n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744;
  wire n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752;
  wire n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760;
  wire n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768;
  wire n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776;
  wire n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784;
  wire n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792;
  wire n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800;
  wire n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808;
  wire n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816;
  wire n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824;
  wire n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832;
  wire n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840;
  wire n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848;
  wire n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856;
  wire n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864;
  wire n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872;
  wire n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880;
  wire n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888;
  wire n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896;
  wire n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904;
  wire n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912;
  wire n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920;
  wire n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928;
  wire n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936;
  wire n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944;
  wire n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952;
  wire n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960;
  wire n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968;
  wire n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976;
  wire n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984;
  wire n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992;
  wire n_3993, n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000;
  wire n_4001, n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008;
  wire n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016;
  wire n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024;
  wire n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032;
  wire n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040;
  wire n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048;
  wire n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056;
  wire n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064;
  wire n_4065, n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072;
  wire n_4073, n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080;
  wire n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088;
  wire n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096;
  wire n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104;
  wire n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112;
  wire n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120;
  wire n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128;
  wire n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136;
  wire n_4137, n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144;
  wire n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152;
  wire n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160;
  wire n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168;
  wire n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176;
  wire n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184;
  wire n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192;
  wire n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200;
  wire n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208;
  wire n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216;
  wire n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224;
  wire n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232;
  wire n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240;
  wire n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248;
  wire n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256;
  wire n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264;
  wire n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272;
  wire n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280;
  wire n_4281, n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288;
  wire n_4289, n_4290, n_4291, n_4292, n_4293, n_4294, n_4295, n_4296;
  wire n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, n_4303, n_4304;
  wire n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312;
  wire n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320;
  wire n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328;
  wire n_4329, n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336;
  wire n_4337, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344;
  wire n_4345, n_4346, n_4347, n_4348, n_4349, n_4350, n_4351, n_4352;
  wire n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360;
  wire n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367, n_4368;
  wire n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376;
  wire n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, n_4384;
  wire n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392;
  wire n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400;
  wire n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408;
  wire n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416;
  wire n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424;
  wire n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432;
  wire n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440;
  wire n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448;
  wire n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456;
  wire n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463, n_4464;
  wire n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472;
  wire n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480;
  wire n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488;
  wire n_4489, n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496;
  wire n_4497, n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504;
  wire n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512;
  wire n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520;
  wire n_4521, n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528;
  wire n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536;
  wire n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544;
  wire n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552;
  wire n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560;
  wire n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568;
  wire n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576;
  wire n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584;
  wire n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592;
  wire n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600;
  wire n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608;
  wire n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616;
  wire n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624;
  wire n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632;
  wire n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640;
  wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648;
  wire n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656;
  wire n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664;
  wire n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672;
  wire n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680;
  wire n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688;
  wire n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696;
  wire n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704;
  wire n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712;
  wire n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720;
  wire n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728;
  wire n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736;
  wire n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744;
  wire n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752;
  wire n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760;
  wire n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768;
  wire n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776;
  wire n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784;
  wire n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792;
  wire n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800;
  wire n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808;
  wire n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816;
  wire n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824;
  wire n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832;
  wire n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840;
  wire n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848;
  wire n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856;
  wire n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864;
  wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872;
  wire n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880;
  wire n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888;
  wire n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896;
  wire n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904;
  wire n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912;
  wire n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920;
  wire n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928;
  wire n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936;
  wire n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944;
  wire n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952;
  wire n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960;
  wire n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968;
  wire n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976;
  wire n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984;
  wire n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992;
  wire n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5000;
  wire n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008;
  wire n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016;
  wire n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024;
  wire n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032;
  wire n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040;
  wire n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048;
  wire n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056;
  wire n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064;
  wire n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072;
  wire n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080;
  wire n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088;
  wire n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096;
  wire n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104;
  wire n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111, n_5112;
  wire n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120;
  wire n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128;
  wire n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136;
  wire n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144;
  wire n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152;
  wire n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160;
  wire n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168;
  wire n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176;
  wire n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184;
  wire n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192;
  wire n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200;
  wire n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208;
  wire n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216;
  wire n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224;
  wire n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232;
  wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
  wire n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248;
  wire n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256;
  wire n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264;
  wire n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272;
  wire n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280;
  wire n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288;
  wire n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296;
  wire n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304;
  wire n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312;
  wire n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320;
  wire n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328;
  wire n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336;
  wire n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344;
  wire n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352;
  wire n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360;
  wire n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368;
  wire n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376;
  wire n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384;
  wire n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392;
  wire n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400;
  wire n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408;
  wire n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416;
  wire n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424;
  wire n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432;
  wire n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440;
  wire n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448;
  wire n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456;
  wire n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464;
  wire n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472;
  wire n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480;
  wire n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488;
  wire n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496;
  wire n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504;
  wire n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512;
  wire n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520;
  wire n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528;
  wire n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536;
  wire n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544;
  wire n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552;
  wire n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560;
  wire n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
  wire n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576;
  wire n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584;
  wire n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592;
  wire n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600;
  wire n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608;
  wire n_5609, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616;
  wire n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624;
  wire n_5625, n_5626, n_5627, n_5628, n_5629, n_5630, n_5631, n_5632;
  wire n_5633, n_5634, n_5635, n_5636, n_5637, n_5638, n_5639, n_5640;
  wire n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5647, n_5648;
  wire n_5649, n_5650, n_5651, n_5652, n_5653, n_5654, n_5655, n_5656;
  wire n_5657, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663, n_5664;
  wire n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672;
  wire n_5673, n_5674, n_5675, n_5676, n_5677, n_5678, n_5679, n_5680;
  wire n_5681, n_5682, n_5683, n_5684, n_5685, n_5686, n_5687, n_5688;
  wire n_5689, n_5690, n_5691, n_5692, n_5693, n_5694, n_5695, n_5696;
  wire n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704;
  wire n_5705, n_5706, n_5707, n_5708, n_5709, n_5710, n_5711, n_5712;
  wire n_5713, n_5714, n_5715, n_5716, n_5717, n_5718, n_5719, n_5720;
  wire n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5727, n_5728;
  wire n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735, n_5736;
  wire n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743, n_5744;
  wire n_5745, n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752;
  wire n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760;
  wire n_5761, n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768;
  wire n_5769, n_5770, n_5771, n_5772, n_5773, n_5774, n_5775, n_5776;
  wire n_5777, n_5778, n_5779, n_5780, n_5781, n_5782, n_5783, n_5784;
  wire n_5785, n_5786, n_5787, n_5788, n_5789, n_5790, n_5791, n_5792;
  wire n_5793, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799, n_5800;
  wire n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5807, n_5808;
  wire n_5809, n_5810, n_5811, n_5812, n_5813, n_5814, n_5815, n_5816;
  wire n_5817, n_5818, n_5819, n_5820, n_5821, n_5822, n_5823, n_5824;
  wire n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831, n_5832;
  wire n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839, n_5840;
  wire n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847, n_5848;
  wire n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5855, n_5856;
  wire n_5857, n_5858, n_5859, n_5860, n_5861, n_5862, n_5863, n_5864;
  wire n_5865, n_5866, n_5867, n_5868, n_5869, n_5870, n_5871, n_5872;
  wire n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880;
  wire n_5881, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888;
  wire n_5889, n_5890, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896;
  wire n_5897, n_5898, n_5899, n_5900, n_5901, n_5902, n_5903, n_5904;
  wire n_5905, n_5906, n_5907, n_5908, n_5909, n_5910, n_5911, n_5912;
  wire n_5913, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919, n_5920;
  wire n_5921, n_5922, n_5923, n_5924, n_5925, n_5926, n_5927, n_5928;
  wire n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935, n_5936;
  wire n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944;
  wire n_5945, n_5946, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952;
  wire n_5953, n_5954, n_5955, n_5956, n_5957, n_5958, n_5959, n_5960;
  wire n_5961, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967, n_5968;
  wire n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975, n_5976;
  wire n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983, n_5984;
  wire n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992;
  wire n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000;
  wire n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008;
  wire n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015, n_6016;
  wire n_6017, n_6018, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024;
  wire n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031, n_6032;
  wire n_6033, n_6034, n_6035, n_6036, n_6037, n_6038, n_6039, n_6040;
  wire n_6041, n_6042, n_6043, n_6044, n_6045, n_6046, n_6047, n_6048;
  wire n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6056;
  wire n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063, n_6064;
  wire n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072;
  wire n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080;
  wire n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087, n_6088;
  wire n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095, n_6096;
  wire n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104;
  wire n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112;
  wire n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120;
  wire n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128;
  wire n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136;
  wire n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144;
  wire n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152;
  wire n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160;
  wire n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168;
  wire n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176;
  wire n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184;
  wire n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192;
  wire n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200;
  wire n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208;
  wire n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216;
  wire n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224;
  wire n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232;
  wire n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240;
  wire n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247, n_6248;
  wire n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256;
  wire n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263, n_6264;
  wire n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271, n_6272;
  wire n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279, n_6280;
  wire n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287, n_6288;
  wire n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295, n_6296;
  wire n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303, n_6304;
  wire n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311, n_6312;
  wire n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319, n_6320;
  wire n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328;
  wire n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336;
  wire n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344;
  wire n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6352;
  wire n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359, n_6360;
  wire n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367, n_6368;
  wire n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376;
  wire n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384;
  wire n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392;
  wire n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400;
  wire n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408;
  wire n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416;
  wire n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424;
  wire n_6425, n_6426, n_6427, n_6428, n_6429, n_6430, n_6431, n_6432;
  wire n_6433, n_6434, n_6435, n_6436, n_6437, n_6438, n_6439, n_6440;
  wire n_6441, n_6442, n_6443, n_6444, n_6445, n_6446, n_6447, n_6448;
  wire n_6449, n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456;
  wire n_6457, n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464;
  wire n_6465, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472;
  wire n_6473, n_6474, n_6475, n_6476, n_6477, n_6478, n_6479, n_6480;
  wire n_6481, n_6482, n_6483, n_6484, n_6485, n_6486, n_6487, n_6488;
  wire n_6489, n_6490, n_6491, n_6492, n_6493, n_6494, n_6495, n_6496;
  wire n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504;
  wire n_6505, n_6506, n_6507, n_6508, n_6509, n_6510, n_6511, n_6512;
  wire n_6513, n_6514, n_6515, n_6516, n_6517, n_6518, n_6519, n_6520;
  wire n_6521, n_6522, n_6523, n_6524, n_6525, n_6526, n_6527, n_6528;
  wire n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536;
  wire n_6537, n_6538, n_6539, n_6540, n_6541, n_6542, n_6543, n_6544;
  wire n_6545, n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6552;
  wire n_6553, n_6554, n_6555, n_6556, n_6557, n_6558, n_6559, n_6560;
  wire n_6561, n_6562, n_6563, n_6564, n_6565, n_6566, n_6567, n_6568;
  wire n_6569, n_6570, n_6571, n_6572, n_6573, n_6574, n_6575, n_6576;
  wire n_6577, n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584;
  wire n_6585, n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592;
  wire n_6593, n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600;
  wire n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608;
  wire n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616;
  wire n_6617, n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624;
  wire n_6625, n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632;
  wire n_6633, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640;
  wire n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648;
  wire n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656;
  wire n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664;
  wire n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672;
  wire n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679, n_6680;
  wire n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688;
  wire n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696;
  wire n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704;
  wire n_6705, n_6706, n_6707, n_6708, n_6709, n_6710, n_6711, n_6712;
  wire n_6713, n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720;
  wire n_6721, n_6722, n_6723, n_6724, n_6725, n_6726, n_6727, n_6728;
  wire n_6729, n_6730, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736;
  wire n_6737, n_6738, n_6739, n_6740, n_6741, n_6742, n_6743, n_6744;
  wire n_6745, n_6746, n_6747, n_6748, n_6749, n_6750, n_6751, n_6752;
  wire n_6753, n_6754, n_6755, n_6756, n_6757, n_6758, n_6759, n_6760;
  wire n_6761, n_6762, n_6763, n_6764, n_6765, n_6766, n_6767, n_6768;
  wire n_6769, n_6770, n_6771, n_6772, n_6773, n_6774, n_6775, n_6776;
  wire n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783, n_6784;
  wire n_6785, n_6786, n_6787, n_6788, n_6789, n_6790, n_6791, n_6792;
  wire n_6793, n_6794, n_6795, n_6796, n_6797, n_6798, n_6799, n_6800;
  wire n_6801, n_6802, n_6803, n_6804, n_6805, n_6806, n_6807, n_6808;
  wire n_6809, n_6810, n_6811, n_6812, n_6813, n_6814, n_6815, n_6816;
  wire n_6817, n_6818, n_6819, n_6820, n_6821, n_6822, n_6823, n_6824;
  wire n_6825, n_6826, n_6827, n_6828, n_6829, n_6830, n_6831, n_6832;
  wire n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6839, n_6840;
  wire n_6841, n_6842, n_6843, n_6844, n_6845, n_6846, n_6847, n_6848;
  wire n_6849, n_6850, n_6851, n_6852, n_6853, n_6854, n_6855, n_6856;
  wire n_6857, n_6858, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864;
  wire n_6865, n_6866, n_6867, n_6868, n_6869, n_6870, n_6871, n_6872;
  wire n_6873, n_6874, n_6875, n_6876, n_6877, n_6878, n_6879, n_6880;
  wire n_6881, n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888;
  wire n_6889, n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896;
  wire n_6897, n_6898, n_6899, n_6900, n_6901, n_6902, n_6903, n_6904;
  wire n_6905, n_6906, n_6907, n_6908, n_6909, n_6910, n_6911, n_6912;
  wire n_6913, n_6914, n_6915, n_6916, n_6917, n_6918, n_6919, n_6920;
  wire n_6921, n_6922, n_6923, n_6924, n_6925, n_6926, n_6927, n_6928;
  wire n_6929, n_6930, n_6931, n_6932, n_6933, n_6934, n_6935, n_6936;
  wire n_6937, n_6938, n_6939, n_6940, n_6941, n_6942, n_6943, n_6944;
  wire n_6945, n_6946, n_6947, n_6948, n_6949, n_6950, n_6951, n_6952;
  wire n_6953, n_6954, n_6955, n_6956, n_6957, n_6958, n_6959, n_6960;
  wire n_6961, n_6962, n_6963, n_6964, n_6965, n_6966, n_6967, n_6968;
  wire n_6969, n_6970, n_6971, n_6972, n_6973, n_6974, n_6975, n_6976;
  wire n_6977, n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984;
  wire n_6985, n_6986, n_6987, n_6988, n_6989, n_6990, n_6991, n_6992;
  wire n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7000;
  wire n_7001, n_7002, n_7003, n_7004, n_7005, n_7006, n_7007, n_7008;
  wire n_7009, n_7010, n_7011, n_7012, n_7013, n_7014, n_7015, n_7016;
  wire n_7017, n_7018, n_7019, n_7020, n_7021, n_7022, n_7023, n_7024;
  wire n_7025, n_7026, n_7027, n_7028, n_7029, n_7030, n_7031, n_7032;
  wire n_7033, n_7034, n_7035, n_7036, n_7037, n_7038, n_7039, n_7040;
  wire n_7041, n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048;
  wire n_7049, n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7056;
  wire n_7057, n_7058, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064;
  wire n_7065, n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072;
  wire n_7073, n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080;
  wire n_7081, n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088;
  wire n_7089, n_7090, n_7091, n_7092, n_7093, n_7094, n_7095, n_7096;
  wire n_7097, n_7098, n_7099, n_7100, n_7101, n_7102, n_7103, n_7104;
  wire n_7105, n_7106, n_7107, n_7108, n_7109, n_7110, n_7111, n_7112;
  wire n_7113, n_7114, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120;
  wire n_7121, n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128;
  wire n_7129, n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136;
  wire n_7137, n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144;
  wire n_7145, n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152;
  wire n_7153, n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7160;
  wire n_7161, n_7162, n_7163, n_7164, n_7165, n_7166, n_7167, n_7168;
  wire n_7169, n_7170, n_7171, n_7172, n_7173, n_7174, n_7175, n_7176;
  wire n_7177, n_7178, n_7179, n_7180, n_7181, n_7182, n_7183, n_7184;
  wire n_7185, n_7186, n_7187, n_7188, n_7189, n_7190, n_7191, n_7192;
  wire n_7193, n_7194, n_7195, n_7196, n_7197, n_7198, n_7199, n_7200;
  wire n_7201, n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208;
  wire n_7209, n_7210, n_7211, n_7212, n_7213, n_7214, n_7215, n_7216;
  wire n_7217, n_7218, n_7219, n_7220, n_7221, n_7222, n_7223, n_7224;
  wire n_7225, n_7226, n_7227, n_7228, n_7229, n_7230, n_7231, n_7232;
  wire n_7233, n_7234, n_7235, n_7236, n_7237, n_7238, n_7239, n_7240;
  wire n_7241, n_7242, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248;
  wire n_7249, n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7256;
  wire n_7257, n_7258, n_7259, n_7260, n_7261, n_7262, n_7263, n_7264;
  wire n_7265, n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272;
  wire n_7273, n_7274, n_7275, n_7276, n_7277, n_7278, n_7279, n_7280;
  wire n_7281, n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288;
  wire n_7289, n_7290, n_7291, n_7292, n_7293, n_7294, n_7295, n_7296;
  wire n_7297, n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304;
  wire n_7305, n_7306, n_7307, n_7308, n_7309, n_7310, n_7311, n_7312;
  wire n_7313, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320;
  wire n_7321, n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328;
  wire n_7329, n_7330, n_7331, n_7332, n_7333, n_7334, n_7335, n_7336;
  wire n_7337, n_7338, n_7339, n_7340, n_7341, n_7342, n_7343, n_7344;
  wire n_7345, n_7346, n_7347, n_7348, n_7349, n_7350, n_7351, n_7352;
  wire n_7353, n_7354, n_7355, n_7356, n_7357, n_7358, n_7359, n_7360;
  wire n_7361, n_7362, n_7363, n_7364, n_7365, n_7366, n_7367, n_7368;
  wire n_7369, n_7370, n_7371, n_7372, n_7373, n_7374, n_7375, n_7376;
  wire n_7377, n_7378, n_7379, n_7380, n_7381, n_7382, n_7383, n_7384;
  wire n_7385, n_7386, n_7387, n_7388, n_7389, n_7390, n_7391, n_7392;
  wire n_7393, n_7394, n_7395, n_7396, n_7397, n_7398, n_7399, n_7400;
  wire n_7401, n_7402, n_7403, n_7404, n_7405, n_7406, n_7407, n_7408;
  wire n_7409, n_7410, n_7411, n_7412, n_7413, n_7414, n_7415, n_7416;
  wire n_7417, n_7418, n_7419, n_7420, n_7421, n_7422, n_7423, n_7424;
  wire n_7425, n_7426, n_7427, n_7428, n_7429, n_7430, n_7431, n_7432;
  wire n_7433, n_7434, n_7435, n_7436, n_7437, n_7438, n_7439, n_7440;
  wire n_7441, n_7442, n_7443, n_7444, n_7445, n_7446, n_7447, n_7448;
  wire n_7449, n_7450, n_7451, n_7452, n_7453, n_7454, n_7455, n_7456;
  wire n_7457, n_7458, n_7459, n_7460, n_7461, n_7462, n_7463, n_7464;
  wire n_7465, n_7466, n_7467, n_7468, n_7469, n_7470, n_7471, n_7472;
  wire n_7473, n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480;
  wire n_7481, n_7482, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488;
  wire n_7489, n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7496;
  wire n_7497, n_7498, n_7499, n_7500, n_7501, n_7502, n_7503, n_7504;
  wire n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_7512;
  wire n_7513, n_7514, n_7515, n_7516, n_7517, n_7518, n_7519, n_7520;
  wire n_7521, n_7522, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528;
  wire n_7529, n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536;
  wire n_7537, n_7538, n_7539, n_7540, n_7541, n_7542, n_7543, n_7544;
  wire n_7545, n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552;
  wire n_7553, n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7560;
  wire n_7561, n_7562, n_7563, n_7564, n_7565, n_7566, n_7567, n_7568;
  wire n_7569, n_7570, n_7571, n_7572, n_7573, n_7574, n_7575, n_7576;
  wire n_7577, n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7584;
  wire n_7585, n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7592;
  wire n_7593, n_7594, n_7595, n_7596, n_7597, n_7598, n_7599, n_7600;
  wire n_7601, n_7602, n_7603, n_7604, n_7605, n_7606, n_7607, n_7608;
  wire n_7609, n_7610, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616;
  wire n_7617, n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624;
  wire n_7625, n_7626, n_7627, n_7628, n_7629, n_7630, n_7631, n_7632;
  wire n_7633, n_7634, n_7635, n_7636, n_7637, n_7638, n_7639, n_7640;
  wire n_7641, n_7642, n_7643, n_7644, n_7645, n_7646, n_7647, n_7648;
  wire n_7649, n_7650, n_7651, n_7652, n_7653, n_7654, n_7655, n_7656;
  wire n_7657, n_7658, n_7659, n_7660, n_7661, n_7662, n_7663, n_7664;
  wire n_7665, n_7666, n_7667, n_7668, n_7669, n_7670, n_7671, n_7672;
  wire n_7673, n_7674, n_7675, n_7676, n_7677, n_7678, n_7679, n_7680;
  wire n_7681, n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688;
  wire n_7689, n_7690, n_7691, n_7692, n_7693, n_7694, n_7695, n_7696;
  wire n_7697, n_7698, n_7699, n_7700, n_7701, n_7702, n_7703, n_7704;
  wire n_7705, n_7706, n_7707, n_7708, n_7709, n_7710, n_7711, n_7712;
  wire n_7713, n_7714, n_7715, n_7716, n_7717, n_7718, n_7719, n_7720;
  wire n_7721, n_7722, n_7723, n_7724, n_7725, n_7726, n_7727, n_7728;
  wire n_7729, n_7730, n_7731, n_7732, n_7733, n_7734, n_7735, n_7736;
  wire n_7737, n_7738, n_7739, n_7740, n_7741, n_7742, n_7743, n_7744;
  wire n_7745, n_7746, n_7747, n_7748, n_7749, n_7750, n_7751, n_7752;
  wire n_7753, n_7754, n_7755, n_7756, n_7757, n_7758, n_7759, n_7760;
  wire n_7761, n_7762, n_7763, n_7764, n_7765, n_7766, n_7767, n_7768;
  wire n_7769, n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776;
  wire n_7777, n_7778, n_7779, n_7780, n_7781, n_7782, n_7783, n_7784;
  wire n_7785, n_7786, n_7787, n_7788, n_7789, n_7790, n_7791, n_7792;
  wire n_7793, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799, n_7800;
  wire n_7801, n_7802, n_7803, n_7804, n_7805, n_7806, n_7807, n_7808;
  wire n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816;
  wire n_7817, n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824;
  wire n_7825, n_7826, n_7827, n_7828, n_7829, n_7830, n_7831, n_7832;
  wire n_7833, n_7834, n_7835, n_7836, n_7837, n_7838, n_7839, n_7840;
  wire n_7841, n_7842, n_7843, n_7844, n_7845, n_7846, n_7847, n_7848;
  wire n_7849, n_7850, n_7851, n_7852, n_7853, n_7854, n_7855, n_7856;
  wire n_7857, n_7858, n_7859, n_7860, n_7861, n_7862, n_7863, n_7864;
  wire n_7865, n_7866, n_7867, n_7868, n_7869, n_7870, n_7871, n_7872;
  wire n_7873, n_7874, n_7875, n_7876, n_7877, n_7878, n_7879, n_7880;
  wire n_7881, n_7882, n_7883, n_7884, n_7885, n_7886, n_7887, n_7888;
  wire n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, n_7895, n_7896;
  wire n_7897, n_7898, n_7899, n_7900, n_7901, n_7902, n_7903, n_7904;
  wire n_7905, n_7906, n_7907, n_7908, n_7909, n_7910, n_7911, n_7912;
  wire n_7913, n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920;
  wire n_7921, n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928;
  wire n_7929, n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936;
  wire n_7937, n_7938, n_7939, n_7940, n_7941, n_7942, n_7943, n_7944;
  wire n_7945, n_7946, n_7947, n_7948, n_7949, n_7950, n_7951, n_7952;
  wire n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960;
  wire n_7961, n_7962, n_7963, n_7964, n_7965, n_7966, n_7967, n_7968;
  wire n_7969, n_7970, n_7971, n_7972, n_7973, n_7974, n_7975, n_7976;
  wire n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983, n_7984;
  wire n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991, n_7992;
  wire n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999, n_8000;
  wire n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007, n_8008;
  wire n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016;
  wire n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024;
  wire n_8025, n_8026, n_8027, n_8028, n_8029, n_8030, n_8031, n_8032;
  wire n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, n_8039, n_8040;
  wire n_8041, n_8042, n_8043, n_8044, n_8045, n_8046, n_8047, n_8048;
  wire n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055, n_8056;
  wire n_8057, n_8058, n_8059, n_8060, n_8061, n_8062, n_8063, n_8064;
  wire n_8065, n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072;
  wire n_8073, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080;
  wire n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088;
  wire n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096;
  wire n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104;
  wire n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112;
  wire n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120;
  wire n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128;
  wire n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136;
  wire n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144;
  wire n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152;
  wire n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160;
  wire n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168;
  wire n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176;
  wire n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184;
  wire n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192;
  wire n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200;
  wire n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208;
  wire n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216;
  wire n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224;
  wire n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232;
  wire n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240;
  wire n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248;
  wire n_8249, n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256;
  wire n_8257, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264;
  wire n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272;
  wire n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280;
  wire n_8281, n_8282, n_8283, n_8284, n_8285, n_8286, n_8287, n_8288;
  wire n_8289, n_8290, n_8291, n_8292, n_8293, n_8294, n_8295, n_8296;
  wire n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304;
  wire n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312;
  wire n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320;
  wire n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328;
  wire n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336;
  wire n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344;
  wire n_8345, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351, n_8352;
  wire n_8353, n_8354, n_8355, n_8356, n_8357, n_8358, n_8359, n_8360;
  wire n_8361, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367, n_8368;
  wire n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376;
  wire n_8377, n_8378, n_8379, n_8380, n_8381, n_8382, n_8383, n_8384;
  wire n_8385, n_8386, n_8387, n_8388, n_8389, n_8390, n_8391, n_8392;
  wire n_8393, n_8394, n_8395, n_8396, n_8397, n_8398, n_8399, n_8400;
  wire n_8401, n_8402, n_8403, n_8404, n_8405, n_8406, n_8407, n_8408;
  wire n_8409, n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416;
  wire n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424;
  wire n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432;
  wire n_8433, n_8434, n_8435, n_8436, n_8437, n_8438, n_8439, n_8440;
  wire n_8441, n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448;
  wire n_8449, n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456;
  wire n_8457, n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464;
  wire n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472;
  wire n_8473, n_8474, n_8475, n_8476, n_8477, n_8478, n_8479, n_8480;
  wire n_8481, n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488;
  wire n_8489, n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496;
  wire n_8497, n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, n_8504;
  wire n_8505, n_8506, n_8507, n_8508, n_8509, n_8510, n_8511, n_8512;
  wire n_8513, n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520;
  wire n_8521, n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528;
  wire n_8529, n_8530, n_8531, n_8532, n_8533, n_8534, n_8535, n_8536;
  wire n_8537, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544;
  wire n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552;
  wire n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560;
  wire n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568;
  wire n_8569, n_8570, n_8571, n_8572, n_8573, n_8574, n_8575, n_8576;
  wire n_8577, n_8578, n_8579, n_8580, n_8581, n_8582, n_8583, n_8584;
  wire n_8585, n_8586, n_8587, n_8588, n_8589, n_8590, n_8591, n_8592;
  wire n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600;
  wire n_8601, n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608;
  wire n_8609, n_8610, n_8611, n_8612, n_8613, n_8614, n_8615, n_8616;
  wire n_8617, n_8618, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624;
  wire n_8625, n_8626, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632;
  wire n_8633, n_8634, n_8635, n_8636, n_8637, n_8638, n_8639, n_8640;
  wire n_8641, n_8642, n_8643, n_8644, n_8645, n_8646, n_8647, n_8648;
  wire n_8649, n_8650, n_8651, n_8652, n_8653, n_8654, n_8655, n_8656;
  wire n_8657, n_8658, n_8659, n_8660, n_8661, n_8662, n_8663, n_8664;
  wire n_8665, n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, n_8672;
  wire n_8673, n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680;
  wire n_8681, n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688;
  wire n_8689, n_8690, n_8691, n_8692, n_8693, n_8694, n_8695, n_8696;
  wire n_8697, n_8698, n_8699, n_8700, n_8701, n_8702, n_8703, n_8704;
  wire n_8705, n_8706, n_8707, n_8708, n_8709, n_8710, n_8711, n_8712;
  wire n_8713, n_8714, n_8715, n_8716, n_8717, n_8718, n_8719, n_8720;
  wire n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727, n_8728;
  wire n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735, n_8736;
  wire n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743, n_8744;
  wire n_8745, n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8752;
  wire n_8753, n_8754, n_8755, n_8756, n_8757, n_8758, n_8759, n_8760;
  wire n_8761, n_8762, n_8763, n_8764, n_8765, n_8766, n_8767, n_8768;
  wire n_8769, n_8770, n_8771, n_8772, n_8773, n_8774, n_8775, n_8776;
  wire n_8777, n_8778, n_8779, n_8780, n_8781, n_8782, n_8783, n_8784;
  wire n_8785, n_8786, n_8787, n_8788, n_8789, n_8790, n_8791, n_8792;
  wire n_8793, n_8794, n_8795, n_8796, n_8797, n_8798, n_8799, n_8800;
  wire n_8801, n_8802, n_8803, n_8804, n_8805, n_8806, n_8807, n_8808;
  wire n_8809, n_8810, n_8811, n_8812, n_8813, n_8814, n_8815, n_8816;
  wire n_8817, n_8818, n_8819, n_8820, n_8821, n_8822, n_8823, n_8824;
  wire n_8825, n_8826, n_8827, n_8828, n_8829, n_8830, n_8831, n_8832;
  wire n_8833, n_8834, n_8835, n_8836, n_8837, n_8838, n_8839, n_8840;
  wire n_8841, n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8848;
  wire n_8849, n_8850, n_8851, n_8852, n_8853, n_8854, n_8855, n_8856;
  wire n_8857, n_8858, n_8859, n_8860, n_8861, n_8862, n_8863, n_8864;
  wire n_8865, n_8866, n_8867, n_8868, n_8869, n_8870, n_8871, n_8872;
  wire n_8873, n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880;
  wire n_8881, n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888;
  wire n_8889, n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896;
  wire n_8897, n_8898, n_8899, n_8900, n_8901, n_8902, n_8903, n_8904;
  wire n_8905, n_8906, n_8907, n_8908, n_8909, n_8910, n_8911, n_8912;
  wire n_8913, n_8914, n_8915, n_8916, n_8917, n_8918, n_8919, n_8920;
  wire n_8921, n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928;
  wire n_8929, n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936;
  wire n_8937, n_8938, n_8939, n_8940, n_8941, n_8942, n_8943, n_8944;
  wire n_8945, n_8946, n_8947, n_8948, n_8949, n_8950, n_8951, n_8952;
  wire n_8953, n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960;
  wire n_8961, n_8962, n_8963, n_8964, n_8965, n_8966, n_8967, n_8968;
  wire n_8969, n_8970, n_8971, n_8972, n_8973, n_8974, n_8975, n_8976;
  wire n_8977, n_8978, n_8979, n_8980, n_8981, n_8982, n_8983, n_8984;
  wire n_8985, n_8986, n_8987, n_8988, n_8989, n_8990, n_8991, n_8992;
  wire n_8993, n_8994, n_8995, n_8996, n_8997, n_8998, n_8999, n_9000;
  wire n_9001, n_9002, n_9003, n_9004, n_9005, n_9006, n_9007, n_9008;
  wire n_9009, n_9010, n_9011, n_9012, n_9013, n_9014, n_9015, n_9016;
  wire n_9017, n_9018, n_9019, n_9020, n_9021, n_9022, n_9023, n_9024;
  wire n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032;
  wire n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040;
  wire n_9041, n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048;
  wire n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056;
  wire n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9064;
  wire n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071, n_9072;
  wire n_9073, n_9074, n_9075, n_9076, n_9077, n_9078, n_9079, n_9080;
  wire n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087, n_9088;
  wire n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095, n_9096;
  wire n_9097, n_9098, n_9099, n_9100, n_9101, n_9102, n_9103, n_9104;
  wire n_9105, n_9106, n_9107, n_9108, n_9109, n_9110, n_9111, n_9112;
  wire n_9113, n_9114, n_9115, n_9116, n_9117, n_9118, n_9119, n_9120;
  wire n_9121, n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128;
  wire n_9129, n_9130, n_9131, n_9132, n_9133, n_9134, n_9135, n_9136;
  wire n_9137, n_9138, n_9139, n_9140, n_9141, n_9142, n_9143, n_9144;
  wire n_9145, n_9146, n_9147, n_9148, n_9149, n_9150, n_9151, n_9152;
  wire n_9153, n_9154, n_9155, n_9156, n_9157, n_9158, n_9159, n_9160;
  wire n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9168;
  wire n_9169, n_9170, n_9171, n_9172, n_9173, n_9174, n_9175, n_9176;
  wire n_9177, n_9178, n_9179, n_9180, n_9181, n_9182, n_9183, n_9184;
  wire n_9185, n_9186, n_9187, n_9188, n_9189, n_9190, n_9191, n_9192;
  wire n_9193, n_9194, n_9195, n_9196, n_9197, n_9198, n_9199, n_9200;
  wire n_9201, n_9202, n_9203, n_9204, n_9205, n_9206, n_9207, n_9208;
  wire n_9209, n_9210, n_9211, n_9212, n_9213, n_9214, n_9215, n_9216;
  wire n_9217, n_9218, n_9219, n_9220, n_9221, n_9222, n_9223, n_9224;
  wire n_9225, n_9226, n_9227, n_9228, n_9229, n_9230, n_9231, n_9232;
  wire n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9239, n_9240;
  wire n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9247, n_9248;
  wire n_9249, n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256;
  wire n_9257, n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264;
  wire n_9265, n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272;
  wire n_9273, n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280;
  wire n_9281, n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288;
  wire n_9289, n_9290, n_9291, n_9292, n_9293, n_9294, n_9295, n_9296;
  wire n_9297, n_9298, n_9299, n_9300, n_9301, n_9302, n_9303, n_9304;
  wire n_9305, n_9306, n_9307, n_9308, n_9309, n_9310, n_9311, n_9312;
  wire n_9313, n_9314, n_9315, n_9316, n_9317, n_9318, n_9319, n_9320;
  wire n_9321, n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9328;
  wire n_9329, n_9330, n_9331, n_9332, n_9333, n_9334, n_9335, n_9336;
  wire n_9337, n_9338, n_9339, n_9340, n_9341, n_9342, n_9343, n_9344;
  wire n_9345, n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352;
  wire n_9353, n_9354, n_9355, n_9356, n_9357, n_9358, n_9359, n_9360;
  wire n_9361, n_9362, n_9363, n_9364, n_9365, n_9366, n_9367, n_9368;
  wire n_9369, n_9370, n_9371, n_9372, n_9373, n_9374, n_9375, n_9376;
  wire n_9377, n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9384;
  wire n_9385, n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, n_9392;
  wire n_9393, n_9394, n_9395, n_9396, n_9397, n_9398, n_9399, n_9400;
  wire n_9401, n_9402, n_9403, n_9404, n_9405, n_9406, n_9407, n_9408;
  wire n_9409, n_9410, n_9411, n_9412, n_9413, n_9414, n_9415, n_9416;
  wire n_9417, n_9418, n_9419, n_9420, n_9421, n_9422, n_9423, n_9424;
  wire n_9425, n_9426, n_9427, n_9428, n_9429, n_9430, n_9431, n_9432;
  wire n_9433, n_9434, n_9435, n_9436, n_9437, n_9438, n_9439, n_9440;
  wire n_9441, n_9442, n_9443, n_9444, n_9445, n_9446, n_9447, n_9448;
  wire n_9449, n_9450, n_9451, n_9452, n_9453, n_9454, n_9455, n_9456;
  wire n_9457, n_9458, n_9459, n_9460, n_9461, n_9462, n_9463, n_9464;
  wire n_9465, n_9466, n_9467, n_9468, n_9469, n_9470, n_9471, n_9472;
  wire n_9473, n_9474, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480;
  wire n_9481, n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488;
  wire n_9489, n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496;
  wire n_9497, n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504;
  wire n_9505, n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512;
  wire n_9513, n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520;
  wire n_9521, n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, n_9528;
  wire n_9529, n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536;
  wire n_9537, n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544;
  wire n_9545, n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552;
  wire n_9553, n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9560;
  wire n_9561, n_9562, n_9563, n_9564, n_9565, n_9566, n_9567, n_9568;
  wire n_9569, n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576;
  wire n_9577, n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584;
  wire n_9585, n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592;
  wire n_9593, n_9594, n_9595, n_9596, n_9597, n_9598, n_9599, n_9600;
  wire n_9601, n_9602, n_9603, n_9604, n_9605, n_9606, n_9607, n_9608;
  wire n_9609, n_9610, n_9611, n_9612, n_9613, n_9614, n_9615, n_9616;
  wire n_9617, n_9618, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624;
  wire n_9625, n_9626, n_9627, n_9628, n_9629, n_9630, n_9631, n_9632;
  wire n_9633, n_9634, n_9635, n_9636, n_9637, n_9638, n_9639, n_9640;
  wire n_9641, n_9642, n_9643, n_9644, n_9645, n_9646, n_9647, n_9648;
  wire n_9649, n_9650, n_9651, n_9652, n_9653, n_9654, n_9655, n_9656;
  wire n_9657, n_9658, n_9659, n_9660, n_9661, n_9662, n_9663, n_9664;
  wire n_9665, n_9666, n_9667, n_9668, n_9669, n_9670, n_9671, n_9672;
  wire n_9673, n_9674, n_9675, n_9676, n_9677, n_9678, n_9679, n_9680;
  wire n_9681, n_9682, n_9683, n_9684, n_9685, n_9686, n_9687, n_9688;
  wire n_9689, n_9690, n_9691, n_9692, n_9693, n_9694, n_9695, n_9696;
  wire n_9697, n_9698, n_9699, n_9700, n_9701, n_9702, n_9703, n_9704;
  wire n_9705, n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712;
  wire n_9713, n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720;
  wire n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728;
  wire n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736;
  wire n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744;
  wire n_9745, n_9746, n_9747, n_9748, n_9749, n_9750, n_9751, n_9752;
  wire n_9753, n_9754, n_9755, n_9756, n_9757, n_9758, n_9759, n_9760;
  wire n_9761, n_9762, n_9763, n_9764, n_9765, n_9766, n_9767, n_9768;
  wire n_9769, n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776;
  wire n_9777, n_9778, n_9779, n_9780, n_9781, n_9782, n_9783, n_9784;
  wire n_9785, n_9786, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792;
  wire n_9793, n_9794, n_9795, n_9796, n_9797, n_9798, n_9799, n_9800;
  wire n_9801, n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808;
  wire n_9809, n_9810, n_9811, n_9812, n_9813, n_9814, n_9815, n_9816;
  wire n_9817, n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824;
  wire n_9825, n_9826, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832;
  wire n_9833, n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840;
  wire n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848;
  wire n_9849, n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856;
  wire n_9857, n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864;
  wire n_9865, n_9866, n_9867, n_9868, n_9869, n_9870, n_9871, n_9872;
  wire n_9873, n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880;
  wire n_9881, n_9882, n_9883, n_9884, n_9885, n_9886, n_9887, n_9888;
  wire n_9889, n_9890, n_9891, n_9892, n_9893, n_9894, n_9895, n_9896;
  wire n_9897, n_9898, n_9899, n_9900, n_9901, n_9902, n_9903, n_9904;
  wire n_9905, n_9906, n_9907, n_9908, n_9909, n_9910, n_9911, n_9912;
  wire n_9913, n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920;
  wire n_9921, n_9922, n_9923, n_9924, n_9925, n_9926, n_9927, n_9928;
  wire n_9929, n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936;
  wire n_9937, n_9938, n_9939, n_9940, n_9941, n_9942, n_9943, n_9944;
  wire n_9945, n_9946, n_9947, n_9948, n_9949, n_9950, n_9951, n_9952;
  wire n_9953, n_9954, n_9955, n_9956, n_9957, n_9958, n_9959, n_9960;
  wire n_9961, n_9962, n_9963, n_9964, n_9965, n_9966, n_9967, n_9968;
  wire n_9969, n_9970, n_9971, n_9972, n_9973, n_9974, n_9975, n_9976;
  wire n_9977, n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984;
  wire n_9985, n_9986, n_9987, n_9988, n_9989, n_9990, n_9991, n_9992;
  wire n_9993, n_9994, n_9995, n_9996, n_9997, n_9998, n_9999, n_10000;
  wire n_10001, n_10002, n_10003, n_10004, n_10005, n_10006, n_10007,
       n_10008;
  wire n_10009, n_10010, n_10011, n_10012, n_10013, n_10014, n_10015,
       n_10016;
  wire n_10017, n_10018, n_10019, n_10020, n_10021, n_10022, n_10023,
       n_10024;
  wire n_10025, n_10026, n_10027, n_10028, n_10029, n_10030, n_10031,
       n_10032;
  wire n_10033, n_10034, n_10035, n_10036, n_10037, n_10038, n_10039,
       n_10040;
  wire n_10041, n_10042, n_10043, n_10044, n_10045, n_10046, n_10047,
       n_10048;
  wire n_10049, n_10050, n_10051, n_10052, n_10053, n_10054, n_10055,
       n_10056;
  wire n_10057, n_10058, n_10059, n_10060, n_10061, n_10062, n_10063,
       n_10064;
  wire n_10065, n_10066, n_10067, n_10068, n_10069, n_10070, n_10071,
       n_10072;
  wire n_10073, n_10074, n_10075, n_10076, n_10077, n_10078, n_10079,
       n_10080;
  wire n_10081, n_10082, n_10083, n_10084, n_10085, n_10086, n_10087,
       n_10088;
  wire n_10089, n_10090, n_10091, n_10092, n_10093, n_10094, n_10095,
       n_10096;
  wire n_10097, n_10098, n_10099, n_10100, n_10101, n_10102, n_10103,
       n_10104;
  wire n_10105, n_10106, n_10107, n_10108, n_10109, n_10110, n_10111,
       n_10112;
  wire n_10113, n_10114, n_10115, n_10116, n_10117, n_10118, n_10119,
       n_10120;
  wire n_10121, n_10122, n_10123, n_10124, n_10125, n_10126, n_10127,
       n_10128;
  wire n_10129, n_10130, n_10131, n_10132, n_10133, n_10134, n_10135,
       n_10136;
  wire n_10137, n_10138, n_10139, n_10140, n_10141, n_10142, n_10143,
       n_10144;
  wire n_10145, n_10146, n_10147, n_10148, n_10149, n_10150, n_10151,
       n_10152;
  wire n_10153, n_10154, n_10155, n_10156, n_10157, n_10158, n_10159,
       n_10160;
  wire n_10161, n_10162, n_10163, n_10164, n_10165, n_10166, n_10167,
       n_10168;
  wire n_10169, n_10170, n_10171, n_10172, n_10173, n_10174, n_10175,
       n_10176;
  wire n_10177, n_10178, n_10179, n_10180, n_10181, n_10182, n_10183,
       n_10184;
  wire n_10185, n_10186, n_10187, n_10188, n_10189, n_10190, n_10191,
       n_10192;
  wire n_10193, n_10194, n_10195, n_10196, n_10197, n_10198, n_10199,
       n_10200;
  wire n_10201, n_10202, n_10203, n_10204, n_10205, n_10206, n_10207,
       n_10208;
  wire n_10209, n_10210, n_10211, n_10212, n_10213, n_10214, n_10215,
       n_10216;
  wire n_10217, n_10218, n_10219, n_10220, n_10221, n_10222, n_10223,
       n_10224;
  wire n_10225, n_10226, n_10227, n_10228, n_10229, n_10230, n_10231,
       n_10232;
  wire n_10233, n_10234, n_10235, n_10236, n_10237, n_10238, n_10239,
       n_10240;
  wire n_10241, n_10242, n_10243, n_10244, n_10245, n_10246, n_10247,
       n_10248;
  wire n_10249, n_10250, n_10251, n_10252, n_10253, n_10254, n_10255,
       n_10256;
  wire n_10257, n_10258, n_10259, n_10260, n_10261, n_10262, n_10263,
       n_10264;
  wire n_10265, n_10266, n_10267, n_10268, n_10269, n_10270, n_10271,
       n_10272;
  wire n_10273, n_10274, n_10275, n_10276, n_10277, n_10278, n_10279,
       n_10280;
  wire n_10281, n_10282, n_10283, n_10284, n_10285, n_10286, n_10287,
       n_10288;
  wire n_10289, n_10290, n_10291, n_10292, n_10293, n_10294, n_10295,
       n_10296;
  wire n_10297, n_10298, n_10299, n_10300, n_10301, n_10302, n_10303,
       n_10304;
  wire n_10305, n_10306, n_10307, n_10308, n_10309, n_10310, n_10311,
       n_10312;
  wire n_10313, n_10314, n_10315, n_10316, n_10317, n_10318, n_10319,
       n_10320;
  wire n_10321, n_10322, n_10323, n_10324, n_10325, n_10326, n_10327,
       n_10328;
  wire n_10329, n_10330, n_10331, n_10332, n_10333, n_10334, n_10335,
       n_10336;
  wire n_10337, n_10338, n_10339, n_10340, n_10341, n_10342, n_10343,
       n_10344;
  wire n_10345, n_10346, n_10347, n_10348, n_10349, n_10350, n_10351,
       n_10352;
  wire n_10353, n_10354, n_10355, n_10356, n_10357, n_10358, n_10359,
       n_10360;
  wire n_10361, n_10362, n_10363, n_10364, n_10365, n_10366, n_10367,
       n_10368;
  wire n_10369, n_10370, n_10371, n_10372, n_10373, n_10374, n_10375,
       n_10376;
  wire n_10377, n_10378, n_10379, n_10380, n_10381, n_10382, n_10383,
       n_10384;
  wire n_10385, n_10386, n_10387, n_10388, n_10389, n_10390, n_10391,
       n_10392;
  wire n_10393, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399,
       n_10400;
  wire n_10401, n_10402, n_10403, n_10404, n_10405, n_10406, n_10407,
       n_10408;
  wire n_10409, n_10410, n_10411, n_10412, n_10413, n_10414, n_10415,
       n_10416;
  wire n_10417, n_10418, n_10419, n_10420, n_10421, n_10422, n_10423,
       n_10424;
  wire n_10425, n_10426, n_10427, n_10428, n_10429, n_10430, n_10431,
       n_10432;
  wire n_10433, n_10434, n_10435, n_10436, n_10437, n_10438, n_10439,
       n_10440;
  wire n_10441, n_10442, n_10443, n_10444, n_10445, n_10446, n_10447,
       n_10448;
  wire n_10449, n_10450, n_10451, n_10452, n_10453, n_10454, n_10455,
       n_10456;
  wire n_10457, n_10458, n_10459, n_10460, n_10461, n_10462, n_10463,
       n_10464;
  wire n_10465, n_10466, n_10467, n_10468, n_10469, n_10470, n_10471,
       n_10472;
  wire n_10473, n_10474, n_10475, n_10476, n_10477, n_10478, n_10479,
       n_10480;
  wire n_10481, n_10482, n_10483, n_10484, n_10485, n_10486, n_10487,
       n_10488;
  wire n_10489, n_10490, n_10491, n_10492, n_10493, n_10494, n_10495,
       n_10496;
  wire n_10497, n_10498, n_10499, n_10500, n_10501, n_10502, n_10503,
       n_10504;
  wire n_10505, n_10506, n_10507, n_10508, n_10509, n_10510, n_10511,
       n_10512;
  wire n_10513, n_10514, n_10515, n_10516, n_10517, n_10518, n_10519,
       n_10520;
  wire n_10521, n_10522, n_10523, n_10524, n_10525, n_10526, n_10527,
       n_10528;
  wire n_10529, n_10530, n_10531, n_10532, n_10533, n_10534, n_10535,
       n_10536;
  wire n_10537, n_10538, n_10539, n_10540, n_10541, n_10542, n_10543,
       n_10544;
  wire n_10545, n_10546, n_10547, n_10548, n_10549, n_10550, n_10551,
       n_10552;
  wire n_10553, n_10554, n_10555, n_10556, n_10557, n_10558, n_10559,
       n_10560;
  wire n_10561, n_10562, n_10563, n_10564, n_10565, n_10566, n_10567,
       n_10568;
  wire n_10569, n_10570, n_10571, n_10572, n_10573, n_10574, n_10575,
       n_10576;
  wire n_10577, n_10578, n_10579, n_10580, n_10581, n_10582, n_10583,
       n_10584;
  wire n_10585, n_10586, n_10587, n_10588, n_10589, n_10590, n_10591,
       n_10592;
  wire n_10593, n_10594, n_10595, n_10596, n_10597, n_10598, n_10599,
       n_10600;
  wire n_10601, n_10602, n_10603, n_10604, n_10605, n_10606, n_10607,
       n_10608;
  wire n_10609, n_10610, n_10611, n_10612, n_10613, n_10614, n_10615,
       n_10616;
  wire n_10617, n_10618, n_10619, n_10620, n_10621, n_10622, n_10623,
       n_10624;
  wire n_10625, n_10626, n_10627, n_10628, n_10629, n_10630, n_10631,
       n_10632;
  wire n_10633, n_10634, n_10635, n_10636, n_10637, n_10638, n_10639,
       n_10640;
  wire n_10641, n_10642, n_10643, n_10644, n_10645, n_10646, n_10647,
       n_10648;
  wire n_10649, n_10650, n_10651, n_10652, n_10653, n_10654, n_10655,
       n_10656;
  wire n_10657, n_10658, n_10659, n_10660, n_10661, n_10662, n_10663,
       n_10664;
  wire n_10665, n_10666, n_10667, n_10668, n_10669, n_10670, n_10671,
       n_10672;
  wire n_10673, n_10674, n_10675, n_10676, n_10677, n_10678, n_10679,
       n_10680;
  wire n_10681, n_10682, n_10683, n_10684, n_10685, n_10686, n_10687,
       n_10688;
  wire n_10689, n_10690, n_10691, n_10692, n_10693, n_10694, n_10695,
       n_10696;
  wire n_10697, n_10698, n_10699, n_10700, n_10701, n_10702, n_10703,
       n_10704;
  wire n_10705, n_10706, n_10707, n_10708, n_10709, n_10710, n_10711,
       n_10712;
  wire n_10713, n_10714, n_10715, n_10716, n_10717, n_10718, n_10719,
       n_10720;
  wire n_10721, n_10722, n_10723, n_10724, n_10725, n_10726, n_10727,
       n_10728;
  wire n_10729, n_10730, n_10731, n_10732, n_10733, n_10734, n_10735,
       n_10736;
  wire n_10737, n_10738, n_10739, n_10740, n_10741, n_10742, n_10743,
       n_10744;
  wire n_10745, n_10746, n_10747, n_10748, n_10749, n_10750, n_10751,
       n_10752;
  wire n_10753, n_10754, n_10755, n_10756, n_10757, n_10758, n_10759,
       n_10760;
  wire n_10761, n_10762, n_10763, n_10764, n_10765, n_10766, n_10767,
       n_10768;
  wire n_10769, n_10770, n_10771, n_10772, n_10773, n_10774, n_10775,
       n_10776;
  wire n_10777, n_10778, n_10779, n_10780, n_10781, n_10782, n_10783,
       n_10784;
  wire n_10785, n_10786, n_10787, n_10788, n_10789, n_10790, n_10791,
       n_10792;
  wire n_10793, n_10794, n_10795, n_10796, n_10797, n_10798, n_10799,
       n_10800;
  wire n_10801, n_10802, n_10803, n_10804, n_10805, n_10806, n_10807,
       n_10808;
  wire n_10809, n_10810, n_10811, n_10812, n_10813, n_10814, n_10815,
       n_10816;
  wire n_10817, n_10818, n_10819, n_10820, n_10821, n_10822, n_10823,
       n_10824;
  wire n_10825, n_10826, n_10827, n_10828, n_10829, n_10830, n_10831,
       n_10832;
  wire n_10833, n_10834, n_10835, n_10836, n_10837, n_10838, n_10839,
       n_10840;
  wire n_10841, n_10842, n_10843, n_10844, n_10845, n_10846, n_10847,
       n_10848;
  wire n_10849, n_10850, n_10851, n_10852, n_10853, n_10854, n_10855,
       n_10856;
  wire n_10857, n_10858, n_10859, n_10860, n_10861, n_10862, n_10863,
       n_10864;
  wire n_10865, n_10866, n_10867, n_10868, n_10869, n_10870, n_10871,
       n_10872;
  wire n_10873, n_10874, n_10875, n_10876, n_10877, n_10878, n_10879,
       n_10880;
  wire n_10881, n_10882, n_10883, n_10884, n_10885, n_10886, n_10887,
       n_10888;
  wire n_10889, n_10890, n_10891, n_10892, n_10893, n_10894, n_10895,
       n_10896;
  wire n_10897, n_10898, n_10899, n_10900, n_10901, n_10902, n_10903,
       n_10904;
  wire n_10905, n_10906, n_10907, n_10908, n_10909, n_10910, n_10911,
       n_10912;
  wire n_10913, n_10914, n_10915, n_10916, n_10917, n_10918, n_10919,
       n_10920;
  wire n_10921, n_10922, n_10923, n_10924, n_10925, n_10926, n_10927,
       n_10928;
  wire n_10929, n_10930, n_10931, n_10932, n_10933, n_10934, n_10935,
       n_10936;
  wire n_10937, n_10938, n_10939, n_10940, n_10941, n_10942, n_10943,
       n_10944;
  wire n_10945, n_10946, n_10947, n_10948, n_10949, n_10950, n_10951,
       n_10952;
  wire n_10953, n_10954, n_10955, n_10956, n_10957, n_10958, n_10959,
       n_10960;
  wire n_10961, n_10962, n_10963, n_10964, n_10965, n_10966, n_10967,
       n_10968;
  wire n_10969, n_10970, n_10971, n_10972, n_10973, n_10974, n_10975,
       n_10976;
  wire n_10977, n_10978, n_10979, n_10980, n_10981, n_10982, n_10983,
       n_10984;
  wire n_10985, n_10986, n_10987, n_10988, n_10989, n_10990, n_10991,
       n_10992;
  wire n_10993, n_10994, n_10995, n_10996, n_10997, n_10998, n_10999,
       n_11000;
  wire n_11001, n_11002, n_11003, n_11004, n_11005, n_11006, n_11007,
       n_11008;
  wire n_11009, n_11010, n_11011, n_11012, n_11013, n_11014, n_11015,
       n_11016;
  wire n_11017, n_11018, n_11019, n_11020, n_11021, n_11022, n_11023,
       n_11024;
  wire n_11025, n_11026, n_11027, n_11028, n_11029, n_11030, n_11031,
       n_11032;
  wire n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, n_11039,
       n_11040;
  wire n_11041, n_11042, n_11043, n_11044, n_11045, n_11046, n_11047,
       n_11048;
  wire n_11049, n_11050, n_11051, n_11052, n_11053, n_11054, n_11055,
       n_11056;
  wire n_11057, n_11058, n_11059, n_11060, n_11061, n_11062, n_11063,
       n_11064;
  wire n_11065, n_11066, n_11067, n_11068, n_11069, n_11070, n_11071,
       n_11072;
  wire n_11073, n_11074, n_11075, n_11076, n_11077, n_11078, n_11079,
       n_11080;
  wire n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087,
       n_11088;
  wire n_11089, n_11090, n_11091, n_11092, n_11093, n_11094, n_11095,
       n_11096;
  wire n_11097, n_11098, n_11099, n_11100, n_11101, n_11102, n_11103,
       n_11104;
  wire n_11105, n_11106, n_11107, n_11108, n_11109, n_11110, n_11111,
       n_11112;
  wire n_11113, n_11114, n_11115, n_11116, n_11117, n_11118, n_11119,
       n_11120;
  wire n_11121, n_11122, n_11123, n_11124, n_11125, n_11126, n_11127,
       n_11128;
  wire n_11129, n_11130, n_11131, n_11132, n_11133, n_11134, n_11135,
       n_11136;
  wire n_11137, n_11138, n_11139, n_11140, n_11141, n_11142, n_11143,
       n_11144;
  wire n_11145, n_11146, n_11147, n_11148, n_11149, n_11150, n_11151,
       n_11152;
  wire n_11153, n_11154, n_11155, n_11156, n_11157, n_11158, n_11159,
       n_11160;
  wire n_11161, n_11162, n_11163, n_11164, n_11165, n_11166, n_11167,
       n_11168;
  wire n_11169, n_11170, n_11171, n_11172, n_11173, n_11174, n_11175,
       n_11176;
  wire n_11177, n_11178, n_11179, n_11180, n_11181, n_11182, n_11183,
       n_11184;
  wire n_11185, n_11186, n_11187, n_11188, n_11189, n_11190, n_11191,
       n_11192;
  wire n_11193, n_11194, n_11195, n_11196, n_11197, n_11198, n_11199,
       n_11200;
  wire n_11201, n_11202, n_11203, n_11204, n_11205, n_11206, n_11207,
       n_11208;
  wire n_11209, n_11210, n_11211, n_11212, n_11213, n_11214, n_11215,
       n_11216;
  wire n_11217, n_11218, n_11219, n_11220, n_11221, n_11222, n_11223,
       n_11224;
  wire n_11225, n_11226, n_11227, n_11228, n_11229, n_11230, n_11231,
       n_11232;
  wire n_11233, n_11234, n_11235, n_11236, n_11237, n_11238, n_11239,
       n_11240;
  wire n_11241, n_11242, n_11243, n_11244, n_11245, n_11246, n_11247,
       n_11248;
  wire n_11249, n_11250, n_11251, n_11252, n_11253, n_11254, n_11255,
       n_11256;
  wire n_11257, n_11258, n_11259, n_11260, n_11261, n_11262, n_11263,
       n_11264;
  wire n_11265, n_11266, n_11267, n_11268, n_11269, n_11270, n_11271,
       n_11272;
  wire n_11273, n_11274, n_11275, n_11276, n_11277, n_11278, n_11279,
       n_11280;
  wire n_11281, n_11282, n_11283, n_11284, n_11285, n_11286, n_11287,
       n_11288;
  wire n_11289, n_11290, n_11291, n_11292, n_11293, n_11294, n_11295,
       n_11296;
  wire n_11297, n_11298, n_11299, n_11300, n_11301, n_11302, n_11303,
       n_11304;
  wire n_11305, n_11306, n_11307, n_11308, n_11309, n_11310, n_11311,
       n_11312;
  wire n_11313, n_11314, n_11315, n_11316, n_11317, n_11318, n_11319,
       n_11320;
  wire n_11321, n_11322, n_11323, n_11324, n_11325, n_11326, n_11327,
       n_11328;
  wire n_11329, n_11330, n_11331, n_11332, n_11333, n_11334, n_11335,
       n_11336;
  wire n_11337, n_11338, n_11339, n_11340, n_11341, n_11342, n_11343,
       n_11344;
  wire n_11345, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351,
       n_11352;
  wire n_11353, n_11354, n_11355, n_11356, n_11357, n_11358, n_11359,
       n_11360;
  wire n_11361, n_11362, n_11363, n_11364, n_11365, n_11366, n_11367,
       n_11368;
  wire n_11369, n_11370, n_11371, n_11372, n_11373, n_11374, n_11375,
       n_11376;
  wire n_11377, n_11378, n_11379, n_11380, n_11381, n_11382, n_11383,
       n_11384;
  wire n_11385, n_11386, n_11387, n_11388, n_11389, n_11390, n_11391,
       n_11392;
  wire n_11393, n_11394, n_11395, n_11396, n_11397, n_11398, n_11399,
       n_11400;
  wire n_11401, n_11402, n_11403, n_11404, n_11405, n_11406, n_11407,
       n_11408;
  wire n_11409, n_11410, n_11411, n_11412, n_11413, n_11414, n_11415,
       n_11416;
  wire n_11417, n_11418, n_11419, n_11420, n_11421, n_11422, n_11423,
       n_11424;
  wire n_11425, n_11426, n_11427, n_11428, n_11429, n_11430, n_11431,
       n_11432;
  wire n_11433, n_11434, n_11435, n_11436, n_11437, n_11438, n_11439,
       n_11440;
  wire n_11441, n_11442, n_11443, n_11444, n_11445, n_11446, n_11447,
       n_11448;
  wire n_11449, n_11450, n_11451, n_11452, n_11453, n_11454, n_11455,
       n_11456;
  wire n_11457, n_11458, n_11459, n_11460, n_11461, n_11462, n_11463,
       n_11464;
  wire n_11465, n_11466, n_11467, n_11468, n_11469, n_11470, n_11471,
       n_11472;
  wire n_11473, n_11474, n_11475, n_11476, n_11477, n_11478, n_11479,
       n_11480;
  wire n_11481, n_11482, n_11483, n_11484, n_11485, n_11486, n_11487,
       n_11488;
  wire n_11489, n_11490, n_11491, n_11492, n_11493, n_11494, n_11495,
       n_11496;
  wire n_11497, n_11498, n_11499, n_11500, n_11501, n_11502, n_11503,
       n_11504;
  wire n_11505, n_11506, n_11507, n_11508, n_11509, n_11510, n_11511,
       n_11512;
  wire n_11513, n_11514, n_11515, n_11516, n_11517, n_11518, n_11519,
       n_11520;
  wire n_11521, n_11522, n_11523, n_11524, n_11525, n_11526, n_11527,
       n_11528;
  wire n_11529, n_11530, n_11531, n_11532, n_11533, n_11534, n_11535,
       n_11536;
  wire n_11537, n_11538, n_11539, n_11540, n_11541, n_11542, n_11543,
       n_11544;
  wire n_11545, n_11546, n_11547, n_11548, n_11549, n_11550, n_11551,
       n_11552;
  wire n_11553, n_11554, n_11555, n_11556, n_11557, n_11558, n_11559,
       n_11560;
  wire n_11561, n_11562, n_11563, n_11564, n_11565, n_11566, n_11567,
       n_11568;
  wire n_11569, n_11570, n_11571, n_11572, n_11573, n_11574, n_11575,
       n_11576;
  wire n_11577, n_11578, n_11579, n_11580, n_11581, n_11582, n_11583,
       n_11584;
  wire n_11585, n_11586, n_11587, n_11588, n_11589, n_11590, n_11591,
       n_11592;
  wire n_11593, n_11594, n_11595, n_11596, n_11597, n_11598, n_11599,
       n_11600;
  wire n_11601, n_11602, n_11603, n_11604, n_11605, n_11606, n_11607,
       n_11608;
  wire n_11609, n_11610, n_11611, n_11612, n_11613, n_11614, n_11615,
       n_11616;
  wire n_11617, n_11618, n_11619, n_11620, n_11621, n_11622, n_11623,
       n_11624;
  wire n_11625, n_11626, n_11627, n_11628, n_11629, n_11630, n_11631,
       n_11632;
  wire n_11633, n_11634, n_11635, n_11636, n_11637, n_11638, n_11639,
       n_11640;
  wire n_11641, n_11642, n_11643, n_11644, n_11645, n_11646, n_11647,
       n_11648;
  wire n_11780, n_11781, n_11782, n_11783, n_11784, n_11785, n_11786,
       n_11787;
  wire n_11788, n_11789, n_11790, n_11791, n_11792, n_11793, n_11794,
       n_11795;
  wire n_11796, n_11797, n_11798, n_11799;
  not g1 (n_3, \req[1] );
  and g2 (n386, \priority[1] , n_3);
  not g3 (n_5, \priority[2] );
  not g4 (n_6, n386);
  and g5 (n387, n_5, n_6);
  not g6 (n_9, \req[2] );
  not g7 (n_10, \req[3] );
  and g8 (n388, n_9, n_10);
  not g9 (n_11, n387);
  and g10 (n389, n_11, n388);
  and g11 (n390, \priority[3] , n_10);
  not g12 (n_14, \priority[4] );
  not g13 (n_15, n390);
  and g14 (n391, n_14, n_15);
  not g15 (n_17, \priority[5] );
  and g16 (n392, n_17, n391);
  not g17 (n_18, n389);
  and g18 (n393, n_18, n392);
  and g19 (n394, n_17, \req[4] );
  not g20 (n_22, \req[5] );
  not g21 (n_23, \req[6] );
  and g22 (n395, n_22, n_23);
  not g23 (n_24, n394);
  and g24 (n396, n_24, n395);
  not g25 (n_25, n393);
  and g26 (n397, n_25, n396);
  and g27 (n398, \priority[6] , n_23);
  not g28 (n_28, \priority[7] );
  not g29 (n_29, n398);
  and g30 (n399, n_28, n_29);
  not g31 (n_31, \priority[8] );
  and g32 (n400, n_31, n399);
  not g33 (n_32, n397);
  and g34 (n401, n_32, n400);
  and g35 (n402, n_31, \req[7] );
  not g36 (n_36, \req[8] );
  not g37 (n_37, \req[9] );
  and g38 (n403, n_36, n_37);
  not g39 (n_38, n402);
  and g40 (n404, n_38, n403);
  not g41 (n_39, n401);
  and g42 (n405, n_39, n404);
  and g43 (n406, \priority[9] , n_37);
  not g44 (n_42, \priority[10] );
  not g45 (n_43, n406);
  and g46 (n407, n_42, n_43);
  not g47 (n_45, \priority[11] );
  and g48 (n408, n_45, n407);
  not g49 (n_46, n405);
  and g50 (n409, n_46, n408);
  and g51 (n410, n_45, \req[10] );
  not g52 (n_50, \req[11] );
  not g53 (n_51, \req[12] );
  and g54 (n411, n_50, n_51);
  not g55 (n_52, n410);
  and g56 (n412, n_52, n411);
  not g57 (n_53, n409);
  and g58 (n413, n_53, n412);
  and g59 (n414, \priority[12] , n_51);
  not g60 (n_56, \priority[13] );
  not g61 (n_57, n414);
  and g62 (n415, n_56, n_57);
  not g63 (n_59, \priority[14] );
  and g64 (n416, n_59, n415);
  not g65 (n_60, n413);
  and g66 (n417, n_60, n416);
  and g67 (n418, n_59, \req[13] );
  not g68 (n_64, \req[14] );
  not g69 (n_65, \req[15] );
  and g70 (n419, n_64, n_65);
  not g71 (n_66, n418);
  and g72 (n420, n_66, n419);
  not g73 (n_67, n417);
  and g74 (n421, n_67, n420);
  and g75 (n422, \priority[15] , n_65);
  not g76 (n_70, \priority[16] );
  not g77 (n_71, n422);
  and g78 (n423, n_70, n_71);
  not g79 (n_73, \priority[17] );
  and g80 (n424, n_73, n423);
  not g81 (n_74, n421);
  and g82 (n425, n_74, n424);
  and g83 (n426, n_73, \req[16] );
  not g84 (n_78, \req[17] );
  not g85 (n_79, \req[18] );
  and g86 (n427, n_78, n_79);
  not g87 (n_80, n426);
  and g88 (n428, n_80, n427);
  not g89 (n_81, n425);
  and g90 (n429, n_81, n428);
  and g91 (n430, \priority[18] , n_79);
  not g92 (n_84, \priority[19] );
  not g93 (n_85, n430);
  and g94 (n431, n_84, n_85);
  not g95 (n_87, \priority[20] );
  and g96 (n432, n_87, n431);
  not g97 (n_88, n429);
  and g98 (n433, n_88, n432);
  and g99 (n434, n_87, \req[19] );
  not g100 (n_92, \req[20] );
  not g101 (n_93, \req[21] );
  and g102 (n435, n_92, n_93);
  not g103 (n_94, n434);
  and g104 (n436, n_94, n435);
  not g105 (n_95, n433);
  and g106 (n437, n_95, n436);
  and g107 (n438, \priority[21] , n_93);
  not g108 (n_98, \priority[22] );
  not g109 (n_99, n438);
  and g110 (n439, n_98, n_99);
  not g111 (n_101, \priority[23] );
  and g112 (n440, n_101, n439);
  not g113 (n_102, n437);
  and g114 (n441, n_102, n440);
  and g115 (n442, n_101, \req[22] );
  not g116 (n_106, \req[23] );
  not g117 (n_107, \req[24] );
  and g118 (n443, n_106, n_107);
  not g119 (n_108, n442);
  and g120 (n444, n_108, n443);
  not g121 (n_109, n441);
  and g122 (n445, n_109, n444);
  and g123 (n446, \priority[24] , n_107);
  not g124 (n_112, \priority[25] );
  not g125 (n_113, n446);
  and g126 (n447, n_112, n_113);
  not g127 (n_115, \priority[26] );
  and g128 (n448, n_115, n447);
  not g129 (n_116, n445);
  and g130 (n449, n_116, n448);
  and g131 (n450, n_115, \req[25] );
  not g132 (n_120, \req[26] );
  not g133 (n_121, \req[27] );
  and g134 (n451, n_120, n_121);
  not g135 (n_122, n450);
  and g136 (n452, n_122, n451);
  not g137 (n_123, n449);
  and g138 (n453, n_123, n452);
  and g139 (n454, \priority[27] , n_121);
  not g140 (n_126, \priority[28] );
  not g141 (n_127, n454);
  and g142 (n455, n_126, n_127);
  not g143 (n_129, \priority[29] );
  and g144 (n456, n_129, n455);
  not g145 (n_130, n453);
  and g146 (n457, n_130, n456);
  and g147 (n458, n_129, \req[28] );
  not g148 (n_134, \req[29] );
  not g149 (n_135, \req[30] );
  and g150 (n459, n_134, n_135);
  not g151 (n_136, n458);
  and g152 (n460, n_136, n459);
  not g153 (n_137, n457);
  and g154 (n461, n_137, n460);
  and g155 (n462, \priority[30] , n_135);
  not g156 (n_140, \priority[31] );
  not g157 (n_141, n462);
  and g158 (n463, n_140, n_141);
  not g159 (n_143, \priority[32] );
  and g160 (n464, n_143, n463);
  not g161 (n_144, n461);
  and g162 (n465, n_144, n464);
  and g163 (n466, n_143, \req[31] );
  not g164 (n_148, \req[32] );
  not g165 (n_149, \req[33] );
  and g166 (n467, n_148, n_149);
  not g167 (n_150, n466);
  and g168 (n468, n_150, n467);
  not g169 (n_151, n465);
  and g170 (n469, n_151, n468);
  and g171 (n470, \priority[33] , n_149);
  not g172 (n_154, \priority[34] );
  not g173 (n_155, n470);
  and g174 (n471, n_154, n_155);
  not g175 (n_157, \priority[35] );
  and g176 (n472, n_157, n471);
  not g177 (n_158, n469);
  and g178 (n473, n_158, n472);
  and g179 (n474, n_157, \req[34] );
  not g180 (n_162, \req[35] );
  not g181 (n_163, \req[36] );
  and g182 (n475, n_162, n_163);
  not g183 (n_164, n474);
  and g184 (n476, n_164, n475);
  not g185 (n_165, n473);
  and g186 (n477, n_165, n476);
  and g187 (n478, \priority[36] , n_163);
  not g188 (n_168, \priority[37] );
  not g189 (n_169, n478);
  and g190 (n479, n_168, n_169);
  not g191 (n_171, \priority[38] );
  and g192 (n480, n_171, n479);
  not g193 (n_172, n477);
  and g194 (n481, n_172, n480);
  and g195 (n482, n_171, \req[37] );
  not g196 (n_176, \req[38] );
  not g197 (n_177, \req[39] );
  and g198 (n483, n_176, n_177);
  not g199 (n_178, n482);
  and g200 (n484, n_178, n483);
  not g201 (n_179, n481);
  and g202 (n485, n_179, n484);
  and g203 (n486, \priority[39] , n_177);
  not g204 (n_182, \priority[40] );
  not g205 (n_183, n486);
  and g206 (n487, n_182, n_183);
  not g207 (n_185, \priority[41] );
  and g208 (n488, n_185, n487);
  not g209 (n_186, n485);
  and g210 (n489, n_186, n488);
  and g211 (n490, n_185, \req[40] );
  not g212 (n_190, \req[41] );
  not g213 (n_191, \req[42] );
  and g214 (n491, n_190, n_191);
  not g215 (n_192, n490);
  and g216 (n492, n_192, n491);
  not g217 (n_193, n489);
  and g218 (n493, n_193, n492);
  and g219 (n494, \priority[42] , n_191);
  not g220 (n_196, \priority[43] );
  not g221 (n_197, n494);
  and g222 (n495, n_196, n_197);
  not g223 (n_199, \priority[44] );
  and g224 (n496, n_199, n495);
  not g225 (n_200, n493);
  and g226 (n497, n_200, n496);
  and g227 (n498, n_199, \req[43] );
  not g228 (n_204, \req[44] );
  not g229 (n_205, \req[45] );
  and g230 (n499, n_204, n_205);
  not g231 (n_206, n498);
  and g232 (n500, n_206, n499);
  not g233 (n_207, n497);
  and g234 (n501, n_207, n500);
  and g235 (n502, \priority[45] , n_205);
  not g236 (n_210, \priority[46] );
  not g237 (n_211, n502);
  and g238 (n503, n_210, n_211);
  not g239 (n_213, \priority[47] );
  and g240 (n504, n_213, n503);
  not g241 (n_214, n501);
  and g242 (n505, n_214, n504);
  and g243 (n506, n_213, \req[46] );
  not g244 (n_218, \req[47] );
  not g245 (n_219, \req[48] );
  and g246 (n507, n_218, n_219);
  not g247 (n_220, n506);
  and g248 (n508, n_220, n507);
  not g249 (n_221, n505);
  and g250 (n509, n_221, n508);
  and g251 (n510, \priority[48] , n_219);
  not g252 (n_224, \priority[49] );
  not g253 (n_225, n510);
  and g254 (n511, n_224, n_225);
  not g255 (n_227, \priority[50] );
  and g256 (n512, n_227, n511);
  not g257 (n_228, n509);
  and g258 (n513, n_228, n512);
  and g259 (n514, n_227, \req[49] );
  not g260 (n_232, \req[50] );
  not g261 (n_233, \req[51] );
  and g262 (n515, n_232, n_233);
  not g263 (n_234, n514);
  and g264 (n516, n_234, n515);
  not g265 (n_235, n513);
  and g266 (n517, n_235, n516);
  and g267 (n518, \priority[51] , n_233);
  not g268 (n_238, \priority[52] );
  not g269 (n_239, n518);
  and g270 (n519, n_238, n_239);
  not g271 (n_241, \priority[53] );
  and g272 (n520, n_241, n519);
  not g273 (n_242, n517);
  and g274 (n521, n_242, n520);
  and g275 (n522, n_241, \req[52] );
  not g276 (n_246, \req[53] );
  not g277 (n_247, \req[54] );
  and g278 (n523, n_246, n_247);
  not g279 (n_248, n522);
  and g280 (n524, n_248, n523);
  not g281 (n_249, n521);
  and g282 (n525, n_249, n524);
  and g283 (n526, \priority[54] , n_247);
  not g284 (n_252, \priority[55] );
  not g285 (n_253, n526);
  and g286 (n527, n_252, n_253);
  not g287 (n_255, \priority[56] );
  and g288 (n528, n_255, n527);
  not g289 (n_256, n525);
  and g290 (n529, n_256, n528);
  and g291 (n530, n_255, \req[55] );
  not g292 (n_260, \req[56] );
  not g293 (n_261, \req[57] );
  and g294 (n531, n_260, n_261);
  not g295 (n_262, n530);
  and g296 (n532, n_262, n531);
  not g297 (n_263, n529);
  and g298 (n533, n_263, n532);
  and g299 (n534, \priority[57] , n_261);
  not g300 (n_266, \priority[58] );
  not g301 (n_267, n534);
  and g302 (n535, n_266, n_267);
  not g303 (n_269, \priority[59] );
  and g304 (n536, n_269, n535);
  not g305 (n_270, n533);
  and g306 (n537, n_270, n536);
  and g307 (n538, n_269, \req[58] );
  not g308 (n_274, \req[59] );
  not g309 (n_275, \req[60] );
  and g310 (n539, n_274, n_275);
  not g311 (n_276, n538);
  and g312 (n540, n_276, n539);
  not g313 (n_277, n537);
  and g314 (n541, n_277, n540);
  and g315 (n542, \priority[60] , n_275);
  not g316 (n_280, \priority[61] );
  not g317 (n_281, n542);
  and g318 (n543, n_280, n_281);
  not g319 (n_283, \priority[62] );
  and g320 (n544, n_283, n543);
  not g321 (n_284, n541);
  and g322 (n545, n_284, n544);
  and g323 (n546, n_283, \req[61] );
  not g324 (n_288, \req[62] );
  not g325 (n_289, \req[63] );
  and g326 (n547, n_288, n_289);
  not g327 (n_290, n546);
  and g328 (n548, n_290, n547);
  not g329 (n_291, n545);
  and g330 (n549, n_291, n548);
  and g331 (n550, \priority[63] , n_289);
  not g332 (n_294, \priority[64] );
  not g333 (n_295, n550);
  and g334 (n551, n_294, n_295);
  not g335 (n_297, \priority[65] );
  and g336 (n552, n_297, n551);
  not g337 (n_298, n549);
  and g338 (n553, n_298, n552);
  and g339 (n554, n_297, \req[64] );
  not g340 (n_302, \req[65] );
  not g341 (n_303, \req[66] );
  and g342 (n555, n_302, n_303);
  not g343 (n_304, n554);
  and g344 (n556, n_304, n555);
  not g345 (n_305, n553);
  and g346 (n557, n_305, n556);
  and g347 (n558, \priority[66] , n_303);
  not g348 (n_308, \priority[67] );
  not g349 (n_309, n558);
  and g350 (n559, n_308, n_309);
  not g351 (n_311, \priority[68] );
  and g352 (n560, n_311, n559);
  not g353 (n_312, n557);
  and g354 (n561, n_312, n560);
  and g355 (n562, n_311, \req[67] );
  not g356 (n_316, \req[68] );
  not g357 (n_317, \req[69] );
  and g358 (n563, n_316, n_317);
  not g359 (n_318, n562);
  and g360 (n564, n_318, n563);
  not g361 (n_319, n561);
  and g362 (n565, n_319, n564);
  and g363 (n566, \priority[69] , n_317);
  not g364 (n_322, \priority[70] );
  not g365 (n_323, n566);
  and g366 (n567, n_322, n_323);
  not g367 (n_325, \priority[71] );
  and g368 (n568, n_325, n567);
  not g369 (n_326, n565);
  and g370 (n569, n_326, n568);
  and g371 (n570, n_325, \req[70] );
  not g372 (n_330, \req[71] );
  not g373 (n_331, \req[72] );
  and g374 (n571, n_330, n_331);
  not g375 (n_332, n570);
  and g376 (n572, n_332, n571);
  not g377 (n_333, n569);
  and g378 (n573, n_333, n572);
  and g379 (n574, \priority[72] , n_331);
  not g380 (n_336, \priority[73] );
  not g381 (n_337, n574);
  and g382 (n575, n_336, n_337);
  not g383 (n_339, \priority[74] );
  and g384 (n576, n_339, n575);
  not g385 (n_340, n573);
  and g386 (n577, n_340, n576);
  and g387 (n578, n_339, \req[73] );
  not g388 (n_344, \req[74] );
  not g389 (n_345, \req[75] );
  and g390 (n579, n_344, n_345);
  not g391 (n_346, n578);
  and g392 (n580, n_346, n579);
  not g393 (n_347, n577);
  and g394 (n581, n_347, n580);
  and g395 (n582, \priority[75] , n_345);
  not g396 (n_350, \priority[76] );
  not g397 (n_351, n582);
  and g398 (n583, n_350, n_351);
  not g399 (n_353, \priority[77] );
  and g400 (n584, n_353, n583);
  not g401 (n_354, n581);
  and g402 (n585, n_354, n584);
  and g403 (n586, n_353, \req[76] );
  not g404 (n_358, \req[77] );
  not g405 (n_359, \req[78] );
  and g406 (n587, n_358, n_359);
  not g407 (n_360, n586);
  and g408 (n588, n_360, n587);
  not g409 (n_361, n585);
  and g410 (n589, n_361, n588);
  and g411 (n590, \priority[78] , n_359);
  not g412 (n_364, \priority[79] );
  not g413 (n_365, n590);
  and g414 (n591, n_364, n_365);
  not g415 (n_367, \priority[80] );
  and g416 (n592, n_367, n591);
  not g417 (n_368, n589);
  and g418 (n593, n_368, n592);
  and g419 (n594, n_367, \req[79] );
  not g420 (n_372, \req[80] );
  not g421 (n_373, \req[81] );
  and g422 (n595, n_372, n_373);
  not g423 (n_374, n594);
  and g424 (n596, n_374, n595);
  not g425 (n_375, n593);
  and g426 (n597, n_375, n596);
  and g427 (n598, \priority[81] , n_373);
  not g428 (n_378, \priority[82] );
  not g429 (n_379, n598);
  and g430 (n599, n_378, n_379);
  not g431 (n_381, \priority[83] );
  and g432 (n600, n_381, n599);
  not g433 (n_382, n597);
  and g434 (n601, n_382, n600);
  and g435 (n602, n_381, \req[82] );
  not g436 (n_386, \req[83] );
  not g437 (n_387, \req[84] );
  and g438 (n603, n_386, n_387);
  not g439 (n_388, n602);
  and g440 (n604, n_388, n603);
  not g441 (n_389, n601);
  and g442 (n605, n_389, n604);
  and g443 (n606, \priority[84] , n_387);
  not g444 (n_392, \priority[85] );
  not g445 (n_393, n606);
  and g446 (n607, n_392, n_393);
  not g447 (n_395, \priority[86] );
  and g448 (n608, n_395, n607);
  not g449 (n_396, n605);
  and g450 (n609, n_396, n608);
  and g451 (n610, n_395, \req[85] );
  not g452 (n_400, \req[86] );
  not g453 (n_401, \req[87] );
  and g454 (n611, n_400, n_401);
  not g455 (n_402, n610);
  and g456 (n612, n_402, n611);
  not g457 (n_403, n609);
  and g458 (n613, n_403, n612);
  and g459 (n614, \priority[87] , n_401);
  not g460 (n_406, \priority[88] );
  not g461 (n_407, n614);
  and g462 (n615, n_406, n_407);
  not g463 (n_409, \priority[89] );
  and g464 (n616, n_409, n615);
  not g465 (n_410, n613);
  and g466 (n617, n_410, n616);
  and g467 (n618, n_409, \req[88] );
  not g468 (n_414, \req[89] );
  not g469 (n_415, \req[90] );
  and g470 (n619, n_414, n_415);
  not g471 (n_416, n618);
  and g472 (n620, n_416, n619);
  not g473 (n_417, n617);
  and g474 (n621, n_417, n620);
  and g475 (n622, \priority[90] , n_415);
  not g476 (n_420, \priority[91] );
  not g477 (n_421, n622);
  and g478 (n623, n_420, n_421);
  not g479 (n_423, \priority[92] );
  and g480 (n624, n_423, n623);
  not g481 (n_424, n621);
  and g482 (n625, n_424, n624);
  and g483 (n626, n_423, \req[91] );
  not g484 (n_428, \req[92] );
  not g485 (n_429, \req[93] );
  and g486 (n627, n_428, n_429);
  not g487 (n_430, n626);
  and g488 (n628, n_430, n627);
  not g489 (n_431, n625);
  and g490 (n629, n_431, n628);
  and g491 (n630, \priority[93] , n_429);
  not g492 (n_434, \priority[94] );
  not g493 (n_435, n630);
  and g494 (n631, n_434, n_435);
  not g495 (n_437, \priority[95] );
  and g496 (n632, n_437, n631);
  not g497 (n_438, n629);
  and g498 (n633, n_438, n632);
  and g499 (n634, n_437, \req[94] );
  not g500 (n_442, \req[95] );
  not g501 (n_443, \req[96] );
  and g502 (n635, n_442, n_443);
  not g503 (n_444, n634);
  and g504 (n636, n_444, n635);
  not g505 (n_445, n633);
  and g506 (n637, n_445, n636);
  and g507 (n638, \priority[96] , n_443);
  not g508 (n_448, \priority[97] );
  not g509 (n_449, n638);
  and g510 (n639, n_448, n_449);
  not g511 (n_451, \priority[98] );
  and g512 (n640, n_451, n639);
  not g513 (n_452, n637);
  and g514 (n641, n_452, n640);
  and g515 (n642, n_451, \req[97] );
  not g516 (n_456, \req[98] );
  not g517 (n_457, \req[99] );
  and g518 (n643, n_456, n_457);
  not g519 (n_458, n642);
  and g520 (n644, n_458, n643);
  not g521 (n_459, n641);
  and g522 (n645, n_459, n644);
  and g523 (n646, \priority[99] , n_457);
  not g524 (n_462, \priority[100] );
  not g525 (n_463, n646);
  and g526 (n647, n_462, n_463);
  not g527 (n_465, \priority[101] );
  and g528 (n648, n_465, n647);
  not g529 (n_466, n645);
  and g530 (n649, n_466, n648);
  and g531 (n650, n_465, \req[100] );
  not g532 (n_470, \req[101] );
  not g533 (n_471, \req[102] );
  and g534 (n651, n_470, n_471);
  not g535 (n_472, n650);
  and g536 (n652, n_472, n651);
  not g537 (n_473, n649);
  and g538 (n653, n_473, n652);
  and g539 (n654, \priority[102] , n_471);
  not g540 (n_476, \priority[103] );
  not g541 (n_477, n654);
  and g542 (n655, n_476, n_477);
  not g543 (n_479, \priority[104] );
  and g544 (n656, n_479, n655);
  not g545 (n_480, n653);
  and g546 (n657, n_480, n656);
  and g547 (n658, n_479, \req[103] );
  not g548 (n_484, \req[104] );
  not g549 (n_485, \req[105] );
  and g550 (n659, n_484, n_485);
  not g551 (n_486, n658);
  and g552 (n660, n_486, n659);
  not g553 (n_487, n657);
  and g554 (n661, n_487, n660);
  and g555 (n662, \priority[105] , n_485);
  not g556 (n_490, \priority[106] );
  not g557 (n_491, n662);
  and g558 (n663, n_490, n_491);
  not g559 (n_493, \priority[107] );
  and g560 (n664, n_493, n663);
  not g561 (n_494, n661);
  and g562 (n665, n_494, n664);
  and g563 (n666, n_493, \req[106] );
  not g564 (n_498, \req[107] );
  not g565 (n_499, \req[108] );
  and g566 (n667, n_498, n_499);
  not g567 (n_500, n666);
  and g568 (n668, n_500, n667);
  not g569 (n_501, n665);
  and g570 (n669, n_501, n668);
  and g571 (n670, \priority[108] , n_499);
  not g572 (n_504, \priority[109] );
  not g573 (n_505, n670);
  and g574 (n671, n_504, n_505);
  not g575 (n_507, \priority[110] );
  and g576 (n672, n_507, n671);
  not g577 (n_508, n669);
  and g578 (n673, n_508, n672);
  and g579 (n674, n_507, \req[109] );
  not g580 (n_512, \req[110] );
  not g581 (n_513, \req[111] );
  and g582 (n675, n_512, n_513);
  not g583 (n_514, n674);
  and g584 (n676, n_514, n675);
  not g585 (n_515, n673);
  and g586 (n677, n_515, n676);
  and g587 (n678, \priority[111] , n_513);
  not g588 (n_518, \priority[112] );
  not g589 (n_519, n678);
  and g590 (n679, n_518, n_519);
  not g591 (n_521, \priority[113] );
  and g592 (n680, n_521, n679);
  not g593 (n_522, n677);
  and g594 (n681, n_522, n680);
  and g595 (n682, n_521, \req[112] );
  not g596 (n_526, \req[113] );
  not g597 (n_527, \req[114] );
  and g598 (n683, n_526, n_527);
  not g599 (n_528, n682);
  and g600 (n684, n_528, n683);
  not g601 (n_529, n681);
  and g602 (n685, n_529, n684);
  and g603 (n686, \priority[114] , n_527);
  not g604 (n_532, \priority[115] );
  not g605 (n_533, n686);
  and g606 (n687, n_532, n_533);
  not g607 (n_535, \priority[116] );
  and g608 (n688, n_535, n687);
  not g609 (n_536, n685);
  and g610 (n689, n_536, n688);
  and g611 (n690, n_535, \req[115] );
  not g612 (n_540, \req[116] );
  not g613 (n_541, \req[117] );
  and g614 (n691, n_540, n_541);
  not g615 (n_542, n690);
  and g616 (n692, n_542, n691);
  not g617 (n_543, n689);
  and g618 (n693, n_543, n692);
  and g619 (n694, \priority[117] , n_541);
  not g620 (n_546, \priority[118] );
  not g621 (n_547, n694);
  and g622 (n695, n_546, n_547);
  not g623 (n_549, \priority[119] );
  and g624 (n696, n_549, n695);
  not g625 (n_550, n693);
  and g626 (n697, n_550, n696);
  and g627 (n698, n_549, \req[118] );
  not g628 (n_554, \req[119] );
  not g629 (n_555, \req[120] );
  and g630 (n699, n_554, n_555);
  not g631 (n_556, n698);
  and g632 (n700, n_556, n699);
  not g633 (n_557, n697);
  and g634 (n701, n_557, n700);
  and g635 (n702, \priority[120] , n_555);
  not g636 (n_560, \priority[121] );
  not g637 (n_561, n702);
  and g638 (n703, n_560, n_561);
  not g639 (n_563, \priority[122] );
  and g640 (n704, n_563, n703);
  not g641 (n_564, n701);
  and g642 (n705, n_564, n704);
  and g643 (n706, n_563, \req[121] );
  not g644 (n_568, \req[122] );
  not g645 (n_569, \req[123] );
  and g646 (n707, n_568, n_569);
  not g647 (n_570, n706);
  and g648 (n708, n_570, n707);
  not g649 (n_571, n705);
  and g650 (n709, n_571, n708);
  and g651 (n710, \priority[123] , n_569);
  not g652 (n_574, \priority[124] );
  not g653 (n_575, n710);
  and g654 (n711, n_574, n_575);
  not g655 (n_577, \priority[125] );
  and g656 (n712, n_577, n711);
  not g657 (n_578, n709);
  and g658 (n713, n_578, n712);
  and g659 (n714, n_577, \req[124] );
  not g660 (n_582, \req[125] );
  not g661 (n_583, \req[126] );
  and g662 (n715, n_582, n_583);
  not g663 (n_584, n714);
  and g664 (n716, n_584, n715);
  not g665 (n_585, n713);
  and g666 (n717, n_585, n716);
  and g667 (n718, \priority[126] , n_583);
  not g668 (n_588, \priority[127] );
  not g669 (n_589, n718);
  and g670 (n719, n_588, n_589);
  not g671 (n_591, \priority[0] );
  and g672 (n720, n_591, n719);
  not g673 (n_592, n717);
  and g674 (n721, n_592, n720);
  and g675 (n722, n_591, \req[127] );
  not g676 (n_595, n722);
  and g677 (n723, \req[0] , n_595);
  not g678 (n_596, n721);
  and g679 (\grant[0] , n_596, n723);
  and g680 (n725, \priority[2] , n_9);
  not g681 (n_597, \priority[3] );
  not g682 (n_598, n725);
  and g683 (n726, n_597, n_598);
  not g684 (n_599, \req[4] );
  and g685 (n727, n_10, n_599);
  not g686 (n_600, n726);
  and g687 (n728, n_600, n727);
  and g688 (n729, \priority[4] , n_599);
  not g689 (n_601, n729);
  and g690 (n730, n_17, n_601);
  not g691 (n_602, \priority[6] );
  and g692 (n731, n_602, n730);
  not g693 (n_603, n728);
  and g694 (n732, n_603, n731);
  and g695 (n733, n_602, \req[5] );
  not g696 (n_604, \req[7] );
  and g697 (n734, n_23, n_604);
  not g698 (n_605, n733);
  and g699 (n735, n_605, n734);
  not g700 (n_606, n732);
  and g701 (n736, n_606, n735);
  and g702 (n737, \priority[7] , n_604);
  not g703 (n_607, n737);
  and g704 (n738, n_31, n_607);
  not g705 (n_608, \priority[9] );
  and g706 (n739, n_608, n738);
  not g707 (n_609, n736);
  and g708 (n740, n_609, n739);
  and g709 (n741, n_608, \req[8] );
  not g710 (n_610, \req[10] );
  and g711 (n742, n_37, n_610);
  not g712 (n_611, n741);
  and g713 (n743, n_611, n742);
  not g714 (n_612, n740);
  and g715 (n744, n_612, n743);
  and g716 (n745, \priority[10] , n_610);
  not g717 (n_613, n745);
  and g718 (n746, n_45, n_613);
  not g719 (n_614, \priority[12] );
  and g720 (n747, n_614, n746);
  not g721 (n_615, n744);
  and g722 (n748, n_615, n747);
  and g723 (n749, n_614, \req[11] );
  not g724 (n_616, \req[13] );
  and g725 (n750, n_51, n_616);
  not g726 (n_617, n749);
  and g727 (n751, n_617, n750);
  not g728 (n_618, n748);
  and g729 (n752, n_618, n751);
  and g730 (n753, \priority[13] , n_616);
  not g731 (n_619, n753);
  and g732 (n754, n_59, n_619);
  not g733 (n_620, \priority[15] );
  and g734 (n755, n_620, n754);
  not g735 (n_621, n752);
  and g736 (n756, n_621, n755);
  and g737 (n757, n_620, \req[14] );
  not g738 (n_622, \req[16] );
  and g739 (n758, n_65, n_622);
  not g740 (n_623, n757);
  and g741 (n759, n_623, n758);
  not g742 (n_624, n756);
  and g743 (n760, n_624, n759);
  and g744 (n761, \priority[16] , n_622);
  not g745 (n_625, n761);
  and g746 (n762, n_73, n_625);
  not g747 (n_626, \priority[18] );
  and g748 (n763, n_626, n762);
  not g749 (n_627, n760);
  and g750 (n764, n_627, n763);
  and g751 (n765, n_626, \req[17] );
  not g752 (n_628, \req[19] );
  and g753 (n766, n_79, n_628);
  not g754 (n_629, n765);
  and g755 (n767, n_629, n766);
  not g756 (n_630, n764);
  and g757 (n768, n_630, n767);
  and g758 (n769, \priority[19] , n_628);
  not g759 (n_631, n769);
  and g760 (n770, n_87, n_631);
  not g761 (n_632, \priority[21] );
  and g762 (n771, n_632, n770);
  not g763 (n_633, n768);
  and g764 (n772, n_633, n771);
  and g765 (n773, n_632, \req[20] );
  not g766 (n_634, \req[22] );
  and g767 (n774, n_93, n_634);
  not g768 (n_635, n773);
  and g769 (n775, n_635, n774);
  not g770 (n_636, n772);
  and g771 (n776, n_636, n775);
  and g772 (n777, \priority[22] , n_634);
  not g773 (n_637, n777);
  and g774 (n778, n_101, n_637);
  not g775 (n_638, \priority[24] );
  and g776 (n779, n_638, n778);
  not g777 (n_639, n776);
  and g778 (n780, n_639, n779);
  and g779 (n781, n_638, \req[23] );
  not g780 (n_640, \req[25] );
  and g781 (n782, n_107, n_640);
  not g782 (n_641, n781);
  and g783 (n783, n_641, n782);
  not g784 (n_642, n780);
  and g785 (n784, n_642, n783);
  and g786 (n785, \priority[25] , n_640);
  not g787 (n_643, n785);
  and g788 (n786, n_115, n_643);
  not g789 (n_644, \priority[27] );
  and g790 (n787, n_644, n786);
  not g791 (n_645, n784);
  and g792 (n788, n_645, n787);
  and g793 (n789, n_644, \req[26] );
  not g794 (n_646, \req[28] );
  and g795 (n790, n_121, n_646);
  not g796 (n_647, n789);
  and g797 (n791, n_647, n790);
  not g798 (n_648, n788);
  and g799 (n792, n_648, n791);
  and g800 (n793, \priority[28] , n_646);
  not g801 (n_649, n793);
  and g802 (n794, n_129, n_649);
  not g803 (n_650, \priority[30] );
  and g804 (n795, n_650, n794);
  not g805 (n_651, n792);
  and g806 (n796, n_651, n795);
  and g807 (n797, n_650, \req[29] );
  not g808 (n_652, \req[31] );
  and g809 (n798, n_135, n_652);
  not g810 (n_653, n797);
  and g811 (n799, n_653, n798);
  not g812 (n_654, n796);
  and g813 (n800, n_654, n799);
  and g814 (n801, \priority[31] , n_652);
  not g815 (n_655, n801);
  and g816 (n802, n_143, n_655);
  not g817 (n_656, \priority[33] );
  and g818 (n803, n_656, n802);
  not g819 (n_657, n800);
  and g820 (n804, n_657, n803);
  and g821 (n805, n_656, \req[32] );
  not g822 (n_658, \req[34] );
  and g823 (n806, n_149, n_658);
  not g824 (n_659, n805);
  and g825 (n807, n_659, n806);
  not g826 (n_660, n804);
  and g827 (n808, n_660, n807);
  and g828 (n809, \priority[34] , n_658);
  not g829 (n_661, n809);
  and g830 (n810, n_157, n_661);
  not g831 (n_662, \priority[36] );
  and g832 (n811, n_662, n810);
  not g833 (n_663, n808);
  and g834 (n812, n_663, n811);
  and g835 (n813, n_662, \req[35] );
  not g836 (n_664, \req[37] );
  and g837 (n814, n_163, n_664);
  not g838 (n_665, n813);
  and g839 (n815, n_665, n814);
  not g840 (n_666, n812);
  and g841 (n816, n_666, n815);
  and g842 (n817, \priority[37] , n_664);
  not g843 (n_667, n817);
  and g844 (n818, n_171, n_667);
  not g845 (n_668, \priority[39] );
  and g846 (n819, n_668, n818);
  not g847 (n_669, n816);
  and g848 (n820, n_669, n819);
  and g849 (n821, n_668, \req[38] );
  not g850 (n_670, \req[40] );
  and g851 (n822, n_177, n_670);
  not g852 (n_671, n821);
  and g853 (n823, n_671, n822);
  not g854 (n_672, n820);
  and g855 (n824, n_672, n823);
  and g856 (n825, \priority[40] , n_670);
  not g857 (n_673, n825);
  and g858 (n826, n_185, n_673);
  not g859 (n_674, \priority[42] );
  and g860 (n827, n_674, n826);
  not g861 (n_675, n824);
  and g862 (n828, n_675, n827);
  and g863 (n829, n_674, \req[41] );
  not g864 (n_676, \req[43] );
  and g865 (n830, n_191, n_676);
  not g866 (n_677, n829);
  and g867 (n831, n_677, n830);
  not g868 (n_678, n828);
  and g869 (n832, n_678, n831);
  and g870 (n833, \priority[43] , n_676);
  not g871 (n_679, n833);
  and g872 (n834, n_199, n_679);
  not g873 (n_680, \priority[45] );
  and g874 (n835, n_680, n834);
  not g875 (n_681, n832);
  and g876 (n836, n_681, n835);
  and g877 (n837, n_680, \req[44] );
  not g878 (n_682, \req[46] );
  and g879 (n838, n_205, n_682);
  not g880 (n_683, n837);
  and g881 (n839, n_683, n838);
  not g882 (n_684, n836);
  and g883 (n840, n_684, n839);
  and g884 (n841, \priority[46] , n_682);
  not g885 (n_685, n841);
  and g886 (n842, n_213, n_685);
  not g887 (n_686, \priority[48] );
  and g888 (n843, n_686, n842);
  not g889 (n_687, n840);
  and g890 (n844, n_687, n843);
  and g891 (n845, n_686, \req[47] );
  not g892 (n_688, \req[49] );
  and g893 (n846, n_219, n_688);
  not g894 (n_689, n845);
  and g895 (n847, n_689, n846);
  not g896 (n_690, n844);
  and g897 (n848, n_690, n847);
  and g898 (n849, \priority[49] , n_688);
  not g899 (n_691, n849);
  and g900 (n850, n_227, n_691);
  not g901 (n_692, \priority[51] );
  and g902 (n851, n_692, n850);
  not g903 (n_693, n848);
  and g904 (n852, n_693, n851);
  and g905 (n853, n_692, \req[50] );
  not g906 (n_694, \req[52] );
  and g907 (n854, n_233, n_694);
  not g908 (n_695, n853);
  and g909 (n855, n_695, n854);
  not g910 (n_696, n852);
  and g911 (n856, n_696, n855);
  and g912 (n857, \priority[52] , n_694);
  not g913 (n_697, n857);
  and g914 (n858, n_241, n_697);
  not g915 (n_698, \priority[54] );
  and g916 (n859, n_698, n858);
  not g917 (n_699, n856);
  and g918 (n860, n_699, n859);
  and g919 (n861, n_698, \req[53] );
  not g920 (n_700, \req[55] );
  and g921 (n862, n_247, n_700);
  not g922 (n_701, n861);
  and g923 (n863, n_701, n862);
  not g924 (n_702, n860);
  and g925 (n864, n_702, n863);
  and g926 (n865, \priority[55] , n_700);
  not g927 (n_703, n865);
  and g928 (n866, n_255, n_703);
  not g929 (n_704, \priority[57] );
  and g930 (n867, n_704, n866);
  not g931 (n_705, n864);
  and g932 (n868, n_705, n867);
  and g933 (n869, n_704, \req[56] );
  not g934 (n_706, \req[58] );
  and g935 (n870, n_261, n_706);
  not g936 (n_707, n869);
  and g937 (n871, n_707, n870);
  not g938 (n_708, n868);
  and g939 (n872, n_708, n871);
  and g940 (n873, \priority[58] , n_706);
  not g941 (n_709, n873);
  and g942 (n874, n_269, n_709);
  not g943 (n_710, \priority[60] );
  and g944 (n875, n_710, n874);
  not g945 (n_711, n872);
  and g946 (n876, n_711, n875);
  and g947 (n877, n_710, \req[59] );
  not g948 (n_712, \req[61] );
  and g949 (n878, n_275, n_712);
  not g950 (n_713, n877);
  and g951 (n879, n_713, n878);
  not g952 (n_714, n876);
  and g953 (n880, n_714, n879);
  and g954 (n881, \priority[61] , n_712);
  not g955 (n_715, n881);
  and g956 (n882, n_283, n_715);
  not g957 (n_716, \priority[63] );
  and g958 (n883, n_716, n882);
  not g959 (n_717, n880);
  and g960 (n884, n_717, n883);
  and g961 (n885, n_716, \req[62] );
  not g962 (n_718, \req[64] );
  and g963 (n886, n_289, n_718);
  not g964 (n_719, n885);
  and g965 (n887, n_719, n886);
  not g966 (n_720, n884);
  and g967 (n888, n_720, n887);
  and g968 (n889, \priority[64] , n_718);
  not g969 (n_721, n889);
  and g970 (n890, n_297, n_721);
  not g971 (n_722, \priority[66] );
  and g972 (n891, n_722, n890);
  not g973 (n_723, n888);
  and g974 (n892, n_723, n891);
  and g975 (n893, n_722, \req[65] );
  not g976 (n_724, \req[67] );
  and g977 (n894, n_303, n_724);
  not g978 (n_725, n893);
  and g979 (n895, n_725, n894);
  not g980 (n_726, n892);
  and g981 (n896, n_726, n895);
  and g982 (n897, \priority[67] , n_724);
  not g983 (n_727, n897);
  and g984 (n898, n_311, n_727);
  not g985 (n_728, \priority[69] );
  and g986 (n899, n_728, n898);
  not g987 (n_729, n896);
  and g988 (n900, n_729, n899);
  and g989 (n901, n_728, \req[68] );
  not g990 (n_730, \req[70] );
  and g991 (n902, n_317, n_730);
  not g992 (n_731, n901);
  and g993 (n903, n_731, n902);
  not g994 (n_732, n900);
  and g995 (n904, n_732, n903);
  and g996 (n905, \priority[70] , n_730);
  not g997 (n_733, n905);
  and g998 (n906, n_325, n_733);
  not g999 (n_734, \priority[72] );
  and g1000 (n907, n_734, n906);
  not g1001 (n_735, n904);
  and g1002 (n908, n_735, n907);
  and g1003 (n909, n_734, \req[71] );
  not g1004 (n_736, \req[73] );
  and g1005 (n910, n_331, n_736);
  not g1006 (n_737, n909);
  and g1007 (n911, n_737, n910);
  not g1008 (n_738, n908);
  and g1009 (n912, n_738, n911);
  and g1010 (n913, \priority[73] , n_736);
  not g1011 (n_739, n913);
  and g1012 (n914, n_339, n_739);
  not g1013 (n_740, \priority[75] );
  and g1014 (n915, n_740, n914);
  not g1015 (n_741, n912);
  and g1016 (n916, n_741, n915);
  and g1017 (n917, n_740, \req[74] );
  not g1018 (n_742, \req[76] );
  and g1019 (n918, n_345, n_742);
  not g1020 (n_743, n917);
  and g1021 (n919, n_743, n918);
  not g1022 (n_744, n916);
  and g1023 (n920, n_744, n919);
  and g1024 (n921, \priority[76] , n_742);
  not g1025 (n_745, n921);
  and g1026 (n922, n_353, n_745);
  not g1027 (n_746, \priority[78] );
  and g1028 (n923, n_746, n922);
  not g1029 (n_747, n920);
  and g1030 (n924, n_747, n923);
  and g1031 (n925, n_746, \req[77] );
  not g1032 (n_748, \req[79] );
  and g1033 (n926, n_359, n_748);
  not g1034 (n_749, n925);
  and g1035 (n927, n_749, n926);
  not g1036 (n_750, n924);
  and g1037 (n928, n_750, n927);
  and g1038 (n929, \priority[79] , n_748);
  not g1039 (n_751, n929);
  and g1040 (n930, n_367, n_751);
  not g1041 (n_752, \priority[81] );
  and g1042 (n931, n_752, n930);
  not g1043 (n_753, n928);
  and g1044 (n932, n_753, n931);
  and g1045 (n933, n_752, \req[80] );
  not g1046 (n_754, \req[82] );
  and g1047 (n934, n_373, n_754);
  not g1048 (n_755, n933);
  and g1049 (n935, n_755, n934);
  not g1050 (n_756, n932);
  and g1051 (n936, n_756, n935);
  and g1052 (n937, \priority[82] , n_754);
  not g1053 (n_757, n937);
  and g1054 (n938, n_381, n_757);
  not g1055 (n_758, \priority[84] );
  and g1056 (n939, n_758, n938);
  not g1057 (n_759, n936);
  and g1058 (n940, n_759, n939);
  and g1059 (n941, n_758, \req[83] );
  not g1060 (n_760, \req[85] );
  and g1061 (n942, n_387, n_760);
  not g1062 (n_761, n941);
  and g1063 (n943, n_761, n942);
  not g1064 (n_762, n940);
  and g1065 (n944, n_762, n943);
  and g1066 (n945, \priority[85] , n_760);
  not g1067 (n_763, n945);
  and g1068 (n946, n_395, n_763);
  not g1069 (n_764, \priority[87] );
  and g1070 (n947, n_764, n946);
  not g1071 (n_765, n944);
  and g1072 (n948, n_765, n947);
  and g1073 (n949, n_764, \req[86] );
  not g1074 (n_766, \req[88] );
  and g1075 (n950, n_401, n_766);
  not g1076 (n_767, n949);
  and g1077 (n951, n_767, n950);
  not g1078 (n_768, n948);
  and g1079 (n952, n_768, n951);
  and g1080 (n953, \priority[88] , n_766);
  not g1081 (n_769, n953);
  and g1082 (n954, n_409, n_769);
  not g1083 (n_770, \priority[90] );
  and g1084 (n955, n_770, n954);
  not g1085 (n_771, n952);
  and g1086 (n956, n_771, n955);
  and g1087 (n957, n_770, \req[89] );
  not g1088 (n_772, \req[91] );
  and g1089 (n958, n_415, n_772);
  not g1090 (n_773, n957);
  and g1091 (n959, n_773, n958);
  not g1092 (n_774, n956);
  and g1093 (n960, n_774, n959);
  and g1094 (n961, \priority[91] , n_772);
  not g1095 (n_775, n961);
  and g1096 (n962, n_423, n_775);
  not g1097 (n_776, \priority[93] );
  and g1098 (n963, n_776, n962);
  not g1099 (n_777, n960);
  and g1100 (n964, n_777, n963);
  and g1101 (n965, n_776, \req[92] );
  not g1102 (n_778, \req[94] );
  and g1103 (n966, n_429, n_778);
  not g1104 (n_779, n965);
  and g1105 (n967, n_779, n966);
  not g1106 (n_780, n964);
  and g1107 (n968, n_780, n967);
  and g1108 (n969, \priority[94] , n_778);
  not g1109 (n_781, n969);
  and g1110 (n970, n_437, n_781);
  not g1111 (n_782, \priority[96] );
  and g1112 (n971, n_782, n970);
  not g1113 (n_783, n968);
  and g1114 (n972, n_783, n971);
  and g1115 (n973, n_782, \req[95] );
  not g1116 (n_784, \req[97] );
  and g1117 (n974, n_443, n_784);
  not g1118 (n_785, n973);
  and g1119 (n975, n_785, n974);
  not g1120 (n_786, n972);
  and g1121 (n976, n_786, n975);
  and g1122 (n977, \priority[97] , n_784);
  not g1123 (n_787, n977);
  and g1124 (n978, n_451, n_787);
  not g1125 (n_788, \priority[99] );
  and g1126 (n979, n_788, n978);
  not g1127 (n_789, n976);
  and g1128 (n980, n_789, n979);
  and g1129 (n981, n_788, \req[98] );
  not g1130 (n_790, \req[100] );
  and g1131 (n982, n_457, n_790);
  not g1132 (n_791, n981);
  and g1133 (n983, n_791, n982);
  not g1134 (n_792, n980);
  and g1135 (n984, n_792, n983);
  and g1136 (n985, \priority[100] , n_790);
  not g1137 (n_793, n985);
  and g1138 (n986, n_465, n_793);
  not g1139 (n_794, \priority[102] );
  and g1140 (n987, n_794, n986);
  not g1141 (n_795, n984);
  and g1142 (n988, n_795, n987);
  and g1143 (n989, n_794, \req[101] );
  not g1144 (n_796, \req[103] );
  and g1145 (n990, n_471, n_796);
  not g1146 (n_797, n989);
  and g1147 (n991, n_797, n990);
  not g1148 (n_798, n988);
  and g1149 (n992, n_798, n991);
  and g1150 (n993, \priority[103] , n_796);
  not g1151 (n_799, n993);
  and g1152 (n994, n_479, n_799);
  not g1153 (n_800, \priority[105] );
  and g1154 (n995, n_800, n994);
  not g1155 (n_801, n992);
  and g1156 (n996, n_801, n995);
  and g1157 (n997, n_800, \req[104] );
  not g1158 (n_802, \req[106] );
  and g1159 (n998, n_485, n_802);
  not g1160 (n_803, n997);
  and g1161 (n999, n_803, n998);
  not g1162 (n_804, n996);
  and g1163 (n1000, n_804, n999);
  and g1164 (n1001, \priority[106] , n_802);
  not g1165 (n_805, n1001);
  and g1166 (n1002, n_493, n_805);
  not g1167 (n_806, \priority[108] );
  and g1168 (n1003, n_806, n1002);
  not g1169 (n_807, n1000);
  and g1170 (n1004, n_807, n1003);
  and g1171 (n1005, n_806, \req[107] );
  not g1172 (n_808, \req[109] );
  and g1173 (n1006, n_499, n_808);
  not g1174 (n_809, n1005);
  and g1175 (n1007, n_809, n1006);
  not g1176 (n_810, n1004);
  and g1177 (n1008, n_810, n1007);
  and g1178 (n1009, \priority[109] , n_808);
  not g1179 (n_811, n1009);
  and g1180 (n1010, n_507, n_811);
  not g1181 (n_812, \priority[111] );
  and g1182 (n1011, n_812, n1010);
  not g1183 (n_813, n1008);
  and g1184 (n1012, n_813, n1011);
  and g1185 (n1013, n_812, \req[110] );
  not g1186 (n_814, \req[112] );
  and g1187 (n1014, n_513, n_814);
  not g1188 (n_815, n1013);
  and g1189 (n1015, n_815, n1014);
  not g1190 (n_816, n1012);
  and g1191 (n1016, n_816, n1015);
  and g1192 (n1017, \priority[112] , n_814);
  not g1193 (n_817, n1017);
  and g1194 (n1018, n_521, n_817);
  not g1195 (n_818, \priority[114] );
  and g1196 (n1019, n_818, n1018);
  not g1197 (n_819, n1016);
  and g1198 (n1020, n_819, n1019);
  and g1199 (n1021, n_818, \req[113] );
  not g1200 (n_820, \req[115] );
  and g1201 (n1022, n_527, n_820);
  not g1202 (n_821, n1021);
  and g1203 (n1023, n_821, n1022);
  not g1204 (n_822, n1020);
  and g1205 (n1024, n_822, n1023);
  and g1206 (n1025, \priority[115] , n_820);
  not g1207 (n_823, n1025);
  and g1208 (n1026, n_535, n_823);
  not g1209 (n_824, \priority[117] );
  and g1210 (n1027, n_824, n1026);
  not g1211 (n_825, n1024);
  and g1212 (n1028, n_825, n1027);
  and g1213 (n1029, n_824, \req[116] );
  not g1214 (n_826, \req[118] );
  and g1215 (n1030, n_541, n_826);
  not g1216 (n_827, n1029);
  and g1217 (n1031, n_827, n1030);
  not g1218 (n_828, n1028);
  and g1219 (n1032, n_828, n1031);
  and g1220 (n1033, \priority[118] , n_826);
  not g1221 (n_829, n1033);
  and g1222 (n1034, n_549, n_829);
  not g1223 (n_830, \priority[120] );
  and g1224 (n1035, n_830, n1034);
  not g1225 (n_831, n1032);
  and g1226 (n1036, n_831, n1035);
  and g1227 (n1037, n_830, \req[119] );
  not g1228 (n_832, \req[121] );
  and g1229 (n1038, n_555, n_832);
  not g1230 (n_833, n1037);
  and g1231 (n1039, n_833, n1038);
  not g1232 (n_834, n1036);
  and g1233 (n1040, n_834, n1039);
  and g1234 (n1041, \priority[121] , n_832);
  not g1235 (n_835, n1041);
  and g1236 (n1042, n_563, n_835);
  not g1237 (n_836, \priority[123] );
  and g1238 (n1043, n_836, n1042);
  not g1239 (n_837, n1040);
  and g1240 (n1044, n_837, n1043);
  and g1241 (n1045, n_836, \req[122] );
  not g1242 (n_838, \req[124] );
  and g1243 (n1046, n_569, n_838);
  not g1244 (n_839, n1045);
  and g1245 (n1047, n_839, n1046);
  not g1246 (n_840, n1044);
  and g1247 (n1048, n_840, n1047);
  and g1248 (n1049, \priority[124] , n_838);
  not g1249 (n_841, n1049);
  and g1250 (n1050, n_577, n_841);
  not g1251 (n_842, \priority[126] );
  and g1252 (n1051, n_842, n1050);
  not g1253 (n_843, n1048);
  and g1254 (n1052, n_843, n1051);
  and g1255 (n1053, n_842, \req[125] );
  not g1256 (n_844, \req[127] );
  and g1257 (n1054, n_583, n_844);
  not g1258 (n_845, n1053);
  and g1259 (n1055, n_845, n1054);
  not g1260 (n_846, n1052);
  and g1261 (n1056, n_846, n1055);
  and g1262 (n1057, \priority[127] , n_844);
  not g1263 (n_847, n1057);
  and g1264 (n1058, n_591, n_847);
  not g1265 (n_848, \priority[1] );
  and g1266 (n1059, n_848, n1058);
  not g1267 (n_849, n1056);
  and g1268 (n1060, n_849, n1059);
  and g1269 (n1061, n_848, \req[0] );
  not g1270 (n_850, n1061);
  and g1271 (n1062, \req[1] , n_850);
  not g1272 (n_851, n1060);
  and g1273 (\grant[1] , n_851, n1062);
  and g1274 (n1064, n_599, n_22);
  not g1275 (n_852, n391);
  and g1276 (n1065, n_852, n1064);
  and g1277 (n1066, \priority[5] , n_22);
  not g1278 (n_853, n1066);
  and g1279 (n1067, n_602, n_853);
  and g1280 (n1068, n_28, n1067);
  not g1281 (n_854, n1065);
  and g1282 (n1069, n_854, n1068);
  and g1283 (n1070, n_28, \req[6] );
  and g1284 (n1071, n_604, n_36);
  not g1285 (n_855, n1070);
  and g1286 (n1072, n_855, n1071);
  not g1287 (n_856, n1069);
  and g1288 (n1073, n_856, n1072);
  and g1289 (n1074, \priority[8] , n_36);
  not g1290 (n_857, n1074);
  and g1291 (n1075, n_608, n_857);
  and g1292 (n1076, n_42, n1075);
  not g1293 (n_858, n1073);
  and g1294 (n1077, n_858, n1076);
  and g1295 (n1078, n_42, \req[9] );
  and g1296 (n1079, n_610, n_50);
  not g1297 (n_859, n1078);
  and g1298 (n1080, n_859, n1079);
  not g1299 (n_860, n1077);
  and g1300 (n1081, n_860, n1080);
  and g1301 (n1082, \priority[11] , n_50);
  not g1302 (n_861, n1082);
  and g1303 (n1083, n_614, n_861);
  and g1304 (n1084, n_56, n1083);
  not g1305 (n_862, n1081);
  and g1306 (n1085, n_862, n1084);
  and g1307 (n1086, n_56, \req[12] );
  and g1308 (n1087, n_616, n_64);
  not g1309 (n_863, n1086);
  and g1310 (n1088, n_863, n1087);
  not g1311 (n_864, n1085);
  and g1312 (n1089, n_864, n1088);
  and g1313 (n1090, \priority[14] , n_64);
  not g1314 (n_865, n1090);
  and g1315 (n1091, n_620, n_865);
  and g1316 (n1092, n_70, n1091);
  not g1317 (n_866, n1089);
  and g1318 (n1093, n_866, n1092);
  and g1319 (n1094, n_70, \req[15] );
  and g1320 (n1095, n_622, n_78);
  not g1321 (n_867, n1094);
  and g1322 (n1096, n_867, n1095);
  not g1323 (n_868, n1093);
  and g1324 (n1097, n_868, n1096);
  and g1325 (n1098, \priority[17] , n_78);
  not g1326 (n_869, n1098);
  and g1327 (n1099, n_626, n_869);
  and g1328 (n1100, n_84, n1099);
  not g1329 (n_870, n1097);
  and g1330 (n1101, n_870, n1100);
  and g1331 (n1102, n_84, \req[18] );
  and g1332 (n1103, n_628, n_92);
  not g1333 (n_871, n1102);
  and g1334 (n1104, n_871, n1103);
  not g1335 (n_872, n1101);
  and g1336 (n1105, n_872, n1104);
  and g1337 (n1106, \priority[20] , n_92);
  not g1338 (n_873, n1106);
  and g1339 (n1107, n_632, n_873);
  and g1340 (n1108, n_98, n1107);
  not g1341 (n_874, n1105);
  and g1342 (n1109, n_874, n1108);
  and g1343 (n1110, n_98, \req[21] );
  and g1344 (n1111, n_634, n_106);
  not g1345 (n_875, n1110);
  and g1346 (n1112, n_875, n1111);
  not g1347 (n_876, n1109);
  and g1348 (n1113, n_876, n1112);
  and g1349 (n1114, \priority[23] , n_106);
  not g1350 (n_877, n1114);
  and g1351 (n1115, n_638, n_877);
  and g1352 (n1116, n_112, n1115);
  not g1353 (n_878, n1113);
  and g1354 (n1117, n_878, n1116);
  and g1355 (n1118, n_112, \req[24] );
  and g1356 (n1119, n_640, n_120);
  not g1357 (n_879, n1118);
  and g1358 (n1120, n_879, n1119);
  not g1359 (n_880, n1117);
  and g1360 (n1121, n_880, n1120);
  and g1361 (n1122, \priority[26] , n_120);
  not g1362 (n_881, n1122);
  and g1363 (n1123, n_644, n_881);
  and g1364 (n1124, n_126, n1123);
  not g1365 (n_882, n1121);
  and g1366 (n1125, n_882, n1124);
  and g1367 (n1126, n_126, \req[27] );
  and g1368 (n1127, n_646, n_134);
  not g1369 (n_883, n1126);
  and g1370 (n1128, n_883, n1127);
  not g1371 (n_884, n1125);
  and g1372 (n1129, n_884, n1128);
  and g1373 (n1130, \priority[29] , n_134);
  not g1374 (n_885, n1130);
  and g1375 (n1131, n_650, n_885);
  and g1376 (n1132, n_140, n1131);
  not g1377 (n_886, n1129);
  and g1378 (n1133, n_886, n1132);
  and g1379 (n1134, n_140, \req[30] );
  and g1380 (n1135, n_652, n_148);
  not g1381 (n_887, n1134);
  and g1382 (n1136, n_887, n1135);
  not g1383 (n_888, n1133);
  and g1384 (n1137, n_888, n1136);
  and g1385 (n1138, \priority[32] , n_148);
  not g1386 (n_889, n1138);
  and g1387 (n1139, n_656, n_889);
  and g1388 (n1140, n_154, n1139);
  not g1389 (n_890, n1137);
  and g1390 (n1141, n_890, n1140);
  and g1391 (n1142, n_154, \req[33] );
  and g1392 (n1143, n_658, n_162);
  not g1393 (n_891, n1142);
  and g1394 (n1144, n_891, n1143);
  not g1395 (n_892, n1141);
  and g1396 (n1145, n_892, n1144);
  and g1397 (n1146, \priority[35] , n_162);
  not g1398 (n_893, n1146);
  and g1399 (n1147, n_662, n_893);
  and g1400 (n1148, n_168, n1147);
  not g1401 (n_894, n1145);
  and g1402 (n1149, n_894, n1148);
  and g1403 (n1150, n_168, \req[36] );
  and g1404 (n1151, n_664, n_176);
  not g1405 (n_895, n1150);
  and g1406 (n1152, n_895, n1151);
  not g1407 (n_896, n1149);
  and g1408 (n1153, n_896, n1152);
  and g1409 (n1154, \priority[38] , n_176);
  not g1410 (n_897, n1154);
  and g1411 (n1155, n_668, n_897);
  and g1412 (n1156, n_182, n1155);
  not g1413 (n_898, n1153);
  and g1414 (n1157, n_898, n1156);
  and g1415 (n1158, n_182, \req[39] );
  and g1416 (n1159, n_670, n_190);
  not g1417 (n_899, n1158);
  and g1418 (n1160, n_899, n1159);
  not g1419 (n_900, n1157);
  and g1420 (n1161, n_900, n1160);
  and g1421 (n1162, \priority[41] , n_190);
  not g1422 (n_901, n1162);
  and g1423 (n1163, n_674, n_901);
  and g1424 (n1164, n_196, n1163);
  not g1425 (n_902, n1161);
  and g1426 (n1165, n_902, n1164);
  and g1427 (n1166, n_196, \req[42] );
  and g1428 (n1167, n_676, n_204);
  not g1429 (n_903, n1166);
  and g1430 (n1168, n_903, n1167);
  not g1431 (n_904, n1165);
  and g1432 (n1169, n_904, n1168);
  and g1433 (n1170, \priority[44] , n_204);
  not g1434 (n_905, n1170);
  and g1435 (n1171, n_680, n_905);
  and g1436 (n1172, n_210, n1171);
  not g1437 (n_906, n1169);
  and g1438 (n1173, n_906, n1172);
  and g1439 (n1174, n_210, \req[45] );
  and g1440 (n1175, n_682, n_218);
  not g1441 (n_907, n1174);
  and g1442 (n1176, n_907, n1175);
  not g1443 (n_908, n1173);
  and g1444 (n1177, n_908, n1176);
  and g1445 (n1178, \priority[47] , n_218);
  not g1446 (n_909, n1178);
  and g1447 (n1179, n_686, n_909);
  and g1448 (n1180, n_224, n1179);
  not g1449 (n_910, n1177);
  and g1450 (n1181, n_910, n1180);
  and g1451 (n1182, n_224, \req[48] );
  and g1452 (n1183, n_688, n_232);
  not g1453 (n_911, n1182);
  and g1454 (n1184, n_911, n1183);
  not g1455 (n_912, n1181);
  and g1456 (n1185, n_912, n1184);
  and g1457 (n1186, \priority[50] , n_232);
  not g1458 (n_913, n1186);
  and g1459 (n1187, n_692, n_913);
  and g1460 (n1188, n_238, n1187);
  not g1461 (n_914, n1185);
  and g1462 (n1189, n_914, n1188);
  and g1463 (n1190, n_238, \req[51] );
  and g1464 (n1191, n_694, n_246);
  not g1465 (n_915, n1190);
  and g1466 (n1192, n_915, n1191);
  not g1467 (n_916, n1189);
  and g1468 (n1193, n_916, n1192);
  and g1469 (n1194, \priority[53] , n_246);
  not g1470 (n_917, n1194);
  and g1471 (n1195, n_698, n_917);
  and g1472 (n1196, n_252, n1195);
  not g1473 (n_918, n1193);
  and g1474 (n1197, n_918, n1196);
  and g1475 (n1198, n_252, \req[54] );
  and g1476 (n1199, n_700, n_260);
  not g1477 (n_919, n1198);
  and g1478 (n1200, n_919, n1199);
  not g1479 (n_920, n1197);
  and g1480 (n1201, n_920, n1200);
  and g1481 (n1202, \priority[56] , n_260);
  not g1482 (n_921, n1202);
  and g1483 (n1203, n_704, n_921);
  and g1484 (n1204, n_266, n1203);
  not g1485 (n_922, n1201);
  and g1486 (n1205, n_922, n1204);
  and g1487 (n1206, n_266, \req[57] );
  and g1488 (n1207, n_706, n_274);
  not g1489 (n_923, n1206);
  and g1490 (n1208, n_923, n1207);
  not g1491 (n_924, n1205);
  and g1492 (n1209, n_924, n1208);
  and g1493 (n1210, \priority[59] , n_274);
  not g1494 (n_925, n1210);
  and g1495 (n1211, n_710, n_925);
  and g1496 (n1212, n_280, n1211);
  not g1497 (n_926, n1209);
  and g1498 (n1213, n_926, n1212);
  and g1499 (n1214, n_280, \req[60] );
  and g1500 (n1215, n_712, n_288);
  not g1501 (n_927, n1214);
  and g1502 (n1216, n_927, n1215);
  not g1503 (n_928, n1213);
  and g1504 (n1217, n_928, n1216);
  and g1505 (n1218, \priority[62] , n_288);
  not g1506 (n_929, n1218);
  and g1507 (n1219, n_716, n_929);
  and g1508 (n1220, n_294, n1219);
  not g1509 (n_930, n1217);
  and g1510 (n1221, n_930, n1220);
  and g1511 (n1222, n_294, \req[63] );
  and g1512 (n1223, n_718, n_302);
  not g1513 (n_931, n1222);
  and g1514 (n1224, n_931, n1223);
  not g1515 (n_932, n1221);
  and g1516 (n1225, n_932, n1224);
  and g1517 (n1226, \priority[65] , n_302);
  not g1518 (n_933, n1226);
  and g1519 (n1227, n_722, n_933);
  and g1520 (n1228, n_308, n1227);
  not g1521 (n_934, n1225);
  and g1522 (n1229, n_934, n1228);
  and g1523 (n1230, n_308, \req[66] );
  and g1524 (n1231, n_724, n_316);
  not g1525 (n_935, n1230);
  and g1526 (n1232, n_935, n1231);
  not g1527 (n_936, n1229);
  and g1528 (n1233, n_936, n1232);
  and g1529 (n1234, \priority[68] , n_316);
  not g1530 (n_937, n1234);
  and g1531 (n1235, n_728, n_937);
  and g1532 (n1236, n_322, n1235);
  not g1533 (n_938, n1233);
  and g1534 (n1237, n_938, n1236);
  and g1535 (n1238, n_322, \req[69] );
  and g1536 (n1239, n_730, n_330);
  not g1537 (n_939, n1238);
  and g1538 (n1240, n_939, n1239);
  not g1539 (n_940, n1237);
  and g1540 (n1241, n_940, n1240);
  and g1541 (n1242, \priority[71] , n_330);
  not g1542 (n_941, n1242);
  and g1543 (n1243, n_734, n_941);
  and g1544 (n1244, n_336, n1243);
  not g1545 (n_942, n1241);
  and g1546 (n1245, n_942, n1244);
  and g1547 (n1246, n_336, \req[72] );
  and g1548 (n1247, n_736, n_344);
  not g1549 (n_943, n1246);
  and g1550 (n1248, n_943, n1247);
  not g1551 (n_944, n1245);
  and g1552 (n1249, n_944, n1248);
  and g1553 (n1250, \priority[74] , n_344);
  not g1554 (n_945, n1250);
  and g1555 (n1251, n_740, n_945);
  and g1556 (n1252, n_350, n1251);
  not g1557 (n_946, n1249);
  and g1558 (n1253, n_946, n1252);
  and g1559 (n1254, n_350, \req[75] );
  and g1560 (n1255, n_742, n_358);
  not g1561 (n_947, n1254);
  and g1562 (n1256, n_947, n1255);
  not g1563 (n_948, n1253);
  and g1564 (n1257, n_948, n1256);
  and g1565 (n1258, \priority[77] , n_358);
  not g1566 (n_949, n1258);
  and g1567 (n1259, n_746, n_949);
  and g1568 (n1260, n_364, n1259);
  not g1569 (n_950, n1257);
  and g1570 (n1261, n_950, n1260);
  and g1571 (n1262, n_364, \req[78] );
  and g1572 (n1263, n_748, n_372);
  not g1573 (n_951, n1262);
  and g1574 (n1264, n_951, n1263);
  not g1575 (n_952, n1261);
  and g1576 (n1265, n_952, n1264);
  and g1577 (n1266, \priority[80] , n_372);
  not g1578 (n_953, n1266);
  and g1579 (n1267, n_752, n_953);
  and g1580 (n1268, n_378, n1267);
  not g1581 (n_954, n1265);
  and g1582 (n1269, n_954, n1268);
  and g1583 (n1270, n_378, \req[81] );
  and g1584 (n1271, n_754, n_386);
  not g1585 (n_955, n1270);
  and g1586 (n1272, n_955, n1271);
  not g1587 (n_956, n1269);
  and g1588 (n1273, n_956, n1272);
  and g1589 (n1274, \priority[83] , n_386);
  not g1590 (n_957, n1274);
  and g1591 (n1275, n_758, n_957);
  and g1592 (n1276, n_392, n1275);
  not g1593 (n_958, n1273);
  and g1594 (n1277, n_958, n1276);
  and g1595 (n1278, n_392, \req[84] );
  and g1596 (n1279, n_760, n_400);
  not g1597 (n_959, n1278);
  and g1598 (n1280, n_959, n1279);
  not g1599 (n_960, n1277);
  and g1600 (n1281, n_960, n1280);
  and g1601 (n1282, \priority[86] , n_400);
  not g1602 (n_961, n1282);
  and g1603 (n1283, n_764, n_961);
  and g1604 (n1284, n_406, n1283);
  not g1605 (n_962, n1281);
  and g1606 (n1285, n_962, n1284);
  and g1607 (n1286, n_406, \req[87] );
  and g1608 (n1287, n_766, n_414);
  not g1609 (n_963, n1286);
  and g1610 (n1288, n_963, n1287);
  not g1611 (n_964, n1285);
  and g1612 (n1289, n_964, n1288);
  and g1613 (n1290, \priority[89] , n_414);
  not g1614 (n_965, n1290);
  and g1615 (n1291, n_770, n_965);
  and g1616 (n1292, n_420, n1291);
  not g1617 (n_966, n1289);
  and g1618 (n1293, n_966, n1292);
  and g1619 (n1294, n_420, \req[90] );
  and g1620 (n1295, n_772, n_428);
  not g1621 (n_967, n1294);
  and g1622 (n1296, n_967, n1295);
  not g1623 (n_968, n1293);
  and g1624 (n1297, n_968, n1296);
  and g1625 (n1298, \priority[92] , n_428);
  not g1626 (n_969, n1298);
  and g1627 (n1299, n_776, n_969);
  and g1628 (n1300, n_434, n1299);
  not g1629 (n_970, n1297);
  and g1630 (n1301, n_970, n1300);
  and g1631 (n1302, n_434, \req[93] );
  and g1632 (n1303, n_778, n_442);
  not g1633 (n_971, n1302);
  and g1634 (n1304, n_971, n1303);
  not g1635 (n_972, n1301);
  and g1636 (n1305, n_972, n1304);
  and g1637 (n1306, \priority[95] , n_442);
  not g1638 (n_973, n1306);
  and g1639 (n1307, n_782, n_973);
  and g1640 (n1308, n_448, n1307);
  not g1641 (n_974, n1305);
  and g1642 (n1309, n_974, n1308);
  and g1643 (n1310, n_448, \req[96] );
  and g1644 (n1311, n_784, n_456);
  not g1645 (n_975, n1310);
  and g1646 (n1312, n_975, n1311);
  not g1647 (n_976, n1309);
  and g1648 (n1313, n_976, n1312);
  and g1649 (n1314, \priority[98] , n_456);
  not g1650 (n_977, n1314);
  and g1651 (n1315, n_788, n_977);
  and g1652 (n1316, n_462, n1315);
  not g1653 (n_978, n1313);
  and g1654 (n1317, n_978, n1316);
  and g1655 (n1318, n_462, \req[99] );
  and g1656 (n1319, n_790, n_470);
  not g1657 (n_979, n1318);
  and g1658 (n1320, n_979, n1319);
  not g1659 (n_980, n1317);
  and g1660 (n1321, n_980, n1320);
  and g1661 (n1322, \priority[101] , n_470);
  not g1662 (n_981, n1322);
  and g1663 (n1323, n_794, n_981);
  and g1664 (n1324, n_476, n1323);
  not g1665 (n_982, n1321);
  and g1666 (n1325, n_982, n1324);
  and g1667 (n1326, n_476, \req[102] );
  and g1668 (n1327, n_796, n_484);
  not g1669 (n_983, n1326);
  and g1670 (n1328, n_983, n1327);
  not g1671 (n_984, n1325);
  and g1672 (n1329, n_984, n1328);
  and g1673 (n1330, \priority[104] , n_484);
  not g1674 (n_985, n1330);
  and g1675 (n1331, n_800, n_985);
  and g1676 (n1332, n_490, n1331);
  not g1677 (n_986, n1329);
  and g1678 (n1333, n_986, n1332);
  and g1679 (n1334, n_490, \req[105] );
  and g1680 (n1335, n_802, n_498);
  not g1681 (n_987, n1334);
  and g1682 (n1336, n_987, n1335);
  not g1683 (n_988, n1333);
  and g1684 (n1337, n_988, n1336);
  and g1685 (n1338, \priority[107] , n_498);
  not g1686 (n_989, n1338);
  and g1687 (n1339, n_806, n_989);
  and g1688 (n1340, n_504, n1339);
  not g1689 (n_990, n1337);
  and g1690 (n1341, n_990, n1340);
  and g1691 (n1342, n_504, \req[108] );
  and g1692 (n1343, n_808, n_512);
  not g1693 (n_991, n1342);
  and g1694 (n1344, n_991, n1343);
  not g1695 (n_992, n1341);
  and g1696 (n1345, n_992, n1344);
  and g1697 (n1346, \priority[110] , n_512);
  not g1698 (n_993, n1346);
  and g1699 (n1347, n_812, n_993);
  and g1700 (n1348, n_518, n1347);
  not g1701 (n_994, n1345);
  and g1702 (n1349, n_994, n1348);
  and g1703 (n1350, n_518, \req[111] );
  and g1704 (n1351, n_814, n_526);
  not g1705 (n_995, n1350);
  and g1706 (n1352, n_995, n1351);
  not g1707 (n_996, n1349);
  and g1708 (n1353, n_996, n1352);
  and g1709 (n1354, \priority[113] , n_526);
  not g1710 (n_997, n1354);
  and g1711 (n1355, n_818, n_997);
  and g1712 (n1356, n_532, n1355);
  not g1713 (n_998, n1353);
  and g1714 (n1357, n_998, n1356);
  and g1715 (n1358, n_532, \req[114] );
  and g1716 (n1359, n_820, n_540);
  not g1717 (n_999, n1358);
  and g1718 (n1360, n_999, n1359);
  not g1719 (n_1000, n1357);
  and g1720 (n1361, n_1000, n1360);
  and g1721 (n1362, \priority[116] , n_540);
  not g1722 (n_1001, n1362);
  and g1723 (n1363, n_824, n_1001);
  and g1724 (n1364, n_546, n1363);
  not g1725 (n_1002, n1361);
  and g1726 (n1365, n_1002, n1364);
  and g1727 (n1366, n_546, \req[117] );
  and g1728 (n1367, n_826, n_554);
  not g1729 (n_1003, n1366);
  and g1730 (n1368, n_1003, n1367);
  not g1731 (n_1004, n1365);
  and g1732 (n1369, n_1004, n1368);
  and g1733 (n1370, \priority[119] , n_554);
  not g1734 (n_1005, n1370);
  and g1735 (n1371, n_830, n_1005);
  and g1736 (n1372, n_560, n1371);
  not g1737 (n_1006, n1369);
  and g1738 (n1373, n_1006, n1372);
  and g1739 (n1374, n_560, \req[120] );
  and g1740 (n1375, n_832, n_568);
  not g1741 (n_1007, n1374);
  and g1742 (n1376, n_1007, n1375);
  not g1743 (n_1008, n1373);
  and g1744 (n1377, n_1008, n1376);
  and g1745 (n1378, \priority[122] , n_568);
  not g1746 (n_1009, n1378);
  and g1747 (n1379, n_836, n_1009);
  and g1748 (n1380, n_574, n1379);
  not g1749 (n_1010, n1377);
  and g1750 (n1381, n_1010, n1380);
  and g1751 (n1382, n_574, \req[123] );
  and g1752 (n1383, n_838, n_582);
  not g1753 (n_1011, n1382);
  and g1754 (n1384, n_1011, n1383);
  not g1755 (n_1012, n1381);
  and g1756 (n1385, n_1012, n1384);
  and g1757 (n1386, \priority[125] , n_582);
  not g1758 (n_1013, n1386);
  and g1759 (n1387, n_842, n_1013);
  and g1760 (n1388, n_588, n1387);
  not g1761 (n_1014, n1385);
  and g1762 (n1389, n_1014, n1388);
  and g1763 (n1390, n_588, \req[126] );
  not g1764 (n_1015, \req[0] );
  and g1765 (n1391, n_1015, n_844);
  not g1766 (n_1016, n1390);
  and g1767 (n1392, n_1016, n1391);
  not g1768 (n_1017, n1389);
  and g1769 (n1393, n_1017, n1392);
  and g1770 (n1394, \priority[0] , n_1015);
  not g1771 (n_1018, n1394);
  and g1772 (n1395, n_848, n_1018);
  and g1773 (n1396, n_5, n1395);
  not g1774 (n_1019, n1393);
  and g1775 (n1397, n_1019, n1396);
  and g1776 (n1398, n_5, \req[1] );
  not g1777 (n_1020, n1398);
  and g1778 (n1399, \req[2] , n_1020);
  not g1779 (n_1021, n1397);
  and g1780 (\grant[2] , n_1021, n1399);
  not g1781 (n_1022, n730);
  and g1782 (n1401, n395, n_1022);
  not g1783 (n_1023, n1401);
  and g1784 (n1402, n400, n_1023);
  not g1785 (n_1024, n1402);
  and g1786 (n1403, n404, n_1024);
  not g1787 (n_1025, n1403);
  and g1788 (n1404, n408, n_1025);
  not g1789 (n_1026, n1404);
  and g1790 (n1405, n412, n_1026);
  not g1791 (n_1027, n1405);
  and g1792 (n1406, n416, n_1027);
  not g1793 (n_1028, n1406);
  and g1794 (n1407, n420, n_1028);
  not g1795 (n_1029, n1407);
  and g1796 (n1408, n424, n_1029);
  not g1797 (n_1030, n1408);
  and g1798 (n1409, n428, n_1030);
  not g1799 (n_1031, n1409);
  and g1800 (n1410, n432, n_1031);
  not g1801 (n_1032, n1410);
  and g1802 (n1411, n436, n_1032);
  not g1803 (n_1033, n1411);
  and g1804 (n1412, n440, n_1033);
  not g1805 (n_1034, n1412);
  and g1806 (n1413, n444, n_1034);
  not g1807 (n_1035, n1413);
  and g1808 (n1414, n448, n_1035);
  not g1809 (n_1036, n1414);
  and g1810 (n1415, n452, n_1036);
  not g1811 (n_1037, n1415);
  and g1812 (n1416, n456, n_1037);
  not g1813 (n_1038, n1416);
  and g1814 (n1417, n460, n_1038);
  not g1815 (n_1039, n1417);
  and g1816 (n1418, n464, n_1039);
  not g1817 (n_1040, n1418);
  and g1818 (n1419, n468, n_1040);
  not g1819 (n_1041, n1419);
  and g1820 (n1420, n472, n_1041);
  not g1821 (n_1042, n1420);
  and g1822 (n1421, n476, n_1042);
  not g1823 (n_1043, n1421);
  and g1824 (n1422, n480, n_1043);
  not g1825 (n_1044, n1422);
  and g1826 (n1423, n484, n_1044);
  not g1827 (n_1045, n1423);
  and g1828 (n1424, n488, n_1045);
  not g1829 (n_1046, n1424);
  and g1830 (n1425, n492, n_1046);
  not g1831 (n_1047, n1425);
  and g1832 (n1426, n496, n_1047);
  not g1833 (n_1048, n1426);
  and g1834 (n1427, n500, n_1048);
  not g1835 (n_1049, n1427);
  and g1836 (n1428, n504, n_1049);
  not g1837 (n_1050, n1428);
  and g1838 (n1429, n508, n_1050);
  not g1839 (n_1051, n1429);
  and g1840 (n1430, n512, n_1051);
  not g1841 (n_1052, n1430);
  and g1842 (n1431, n516, n_1052);
  not g1843 (n_1053, n1431);
  and g1844 (n1432, n520, n_1053);
  not g1845 (n_1054, n1432);
  and g1846 (n1433, n524, n_1054);
  not g1847 (n_1055, n1433);
  and g1848 (n1434, n528, n_1055);
  not g1849 (n_1056, n1434);
  and g1850 (n1435, n532, n_1056);
  not g1851 (n_1057, n1435);
  and g1852 (n1436, n536, n_1057);
  not g1853 (n_1058, n1436);
  and g1854 (n1437, n540, n_1058);
  not g1855 (n_1059, n1437);
  and g1856 (n1438, n544, n_1059);
  not g1857 (n_1060, n1438);
  and g1858 (n1439, n548, n_1060);
  not g1859 (n_1061, n1439);
  and g1860 (n1440, n552, n_1061);
  not g1861 (n_1062, n1440);
  and g1862 (n1441, n556, n_1062);
  not g1863 (n_1063, n1441);
  and g1864 (n1442, n560, n_1063);
  not g1865 (n_1064, n1442);
  and g1866 (n1443, n564, n_1064);
  not g1867 (n_1065, n1443);
  and g1868 (n1444, n568, n_1065);
  not g1869 (n_1066, n1444);
  and g1870 (n1445, n572, n_1066);
  not g1871 (n_1067, n1445);
  and g1872 (n1446, n576, n_1067);
  not g1873 (n_1068, n1446);
  and g1874 (n1447, n580, n_1068);
  not g1875 (n_1069, n1447);
  and g1876 (n1448, n584, n_1069);
  not g1877 (n_1070, n1448);
  and g1878 (n1449, n588, n_1070);
  not g1879 (n_1071, n1449);
  and g1880 (n1450, n592, n_1071);
  not g1881 (n_1072, n1450);
  and g1882 (n1451, n596, n_1072);
  not g1883 (n_1073, n1451);
  and g1884 (n1452, n600, n_1073);
  not g1885 (n_1074, n1452);
  and g1886 (n1453, n604, n_1074);
  not g1887 (n_1075, n1453);
  and g1888 (n1454, n608, n_1075);
  not g1889 (n_1076, n1454);
  and g1890 (n1455, n612, n_1076);
  not g1891 (n_1077, n1455);
  and g1892 (n1456, n616, n_1077);
  not g1893 (n_1078, n1456);
  and g1894 (n1457, n620, n_1078);
  not g1895 (n_1079, n1457);
  and g1896 (n1458, n624, n_1079);
  not g1897 (n_1080, n1458);
  and g1898 (n1459, n628, n_1080);
  not g1899 (n_1081, n1459);
  and g1900 (n1460, n632, n_1081);
  not g1901 (n_1082, n1460);
  and g1902 (n1461, n636, n_1082);
  not g1903 (n_1083, n1461);
  and g1904 (n1462, n640, n_1083);
  not g1905 (n_1084, n1462);
  and g1906 (n1463, n644, n_1084);
  not g1907 (n_1085, n1463);
  and g1908 (n1464, n648, n_1085);
  not g1909 (n_1086, n1464);
  and g1910 (n1465, n652, n_1086);
  not g1911 (n_1087, n1465);
  and g1912 (n1466, n656, n_1087);
  not g1913 (n_1088, n1466);
  and g1914 (n1467, n660, n_1088);
  not g1915 (n_1089, n1467);
  and g1916 (n1468, n664, n_1089);
  not g1917 (n_1090, n1468);
  and g1918 (n1469, n668, n_1090);
  not g1919 (n_1091, n1469);
  and g1920 (n1470, n672, n_1091);
  not g1921 (n_1092, n1470);
  and g1922 (n1471, n676, n_1092);
  not g1923 (n_1093, n1471);
  and g1924 (n1472, n680, n_1093);
  not g1925 (n_1094, n1472);
  and g1926 (n1473, n684, n_1094);
  not g1927 (n_1095, n1473);
  and g1928 (n1474, n688, n_1095);
  not g1929 (n_1096, n1474);
  and g1930 (n1475, n692, n_1096);
  not g1931 (n_1097, n1475);
  and g1932 (n1476, n696, n_1097);
  not g1933 (n_1098, n1476);
  and g1934 (n1477, n700, n_1098);
  not g1935 (n_1099, n1477);
  and g1936 (n1478, n704, n_1099);
  not g1937 (n_1100, n1478);
  and g1938 (n1479, n708, n_1100);
  not g1939 (n_1101, n1479);
  and g1940 (n1480, n712, n_1101);
  not g1941 (n_1102, n1480);
  and g1942 (n1481, n716, n_1102);
  not g1943 (n_1103, n1481);
  and g1944 (n1482, n720, n_1103);
  and g1945 (n1483, n_1015, n_3);
  and g1946 (n1484, n_595, n1483);
  not g1947 (n_1104, n1482);
  and g1948 (n1485, n_1104, n1484);
  and g1949 (n1486, n_597, n387);
  not g1950 (n_1105, n1485);
  and g1951 (n1487, n_1105, n1486);
  and g1952 (n1488, n_597, \req[2] );
  not g1953 (n_1106, n1488);
  and g1954 (n1489, \req[3] , n_1106);
  not g1955 (n_1107, n1487);
  and g1956 (\grant[3] , n_1107, n1489);
  not g1957 (n_1108, n1067);
  and g1958 (n1491, n734, n_1108);
  not g1959 (n_1109, n1491);
  and g1960 (n1492, n739, n_1109);
  not g1961 (n_1110, n1492);
  and g1962 (n1493, n743, n_1110);
  not g1963 (n_1111, n1493);
  and g1964 (n1494, n747, n_1111);
  not g1965 (n_1112, n1494);
  and g1966 (n1495, n751, n_1112);
  not g1967 (n_1113, n1495);
  and g1968 (n1496, n755, n_1113);
  not g1969 (n_1114, n1496);
  and g1970 (n1497, n759, n_1114);
  not g1971 (n_1115, n1497);
  and g1972 (n1498, n763, n_1115);
  not g1973 (n_1116, n1498);
  and g1974 (n1499, n767, n_1116);
  not g1975 (n_1117, n1499);
  and g1976 (n1500, n771, n_1117);
  not g1977 (n_1118, n1500);
  and g1978 (n1501, n775, n_1118);
  not g1979 (n_1119, n1501);
  and g1980 (n1502, n779, n_1119);
  not g1981 (n_1120, n1502);
  and g1982 (n1503, n783, n_1120);
  not g1983 (n_1121, n1503);
  and g1984 (n1504, n787, n_1121);
  not g1985 (n_1122, n1504);
  and g1986 (n1505, n791, n_1122);
  not g1987 (n_1123, n1505);
  and g1988 (n1506, n795, n_1123);
  not g1989 (n_1124, n1506);
  and g1990 (n1507, n799, n_1124);
  not g1991 (n_1125, n1507);
  and g1992 (n1508, n803, n_1125);
  not g1993 (n_1126, n1508);
  and g1994 (n1509, n807, n_1126);
  not g1995 (n_1127, n1509);
  and g1996 (n1510, n811, n_1127);
  not g1997 (n_1128, n1510);
  and g1998 (n1511, n815, n_1128);
  not g1999 (n_1129, n1511);
  and g2000 (n1512, n819, n_1129);
  not g2001 (n_1130, n1512);
  and g2002 (n1513, n823, n_1130);
  not g2003 (n_1131, n1513);
  and g2004 (n1514, n827, n_1131);
  not g2005 (n_1132, n1514);
  and g2006 (n1515, n831, n_1132);
  not g2007 (n_1133, n1515);
  and g2008 (n1516, n835, n_1133);
  not g2009 (n_1134, n1516);
  and g2010 (n1517, n839, n_1134);
  not g2011 (n_1135, n1517);
  and g2012 (n1518, n843, n_1135);
  not g2013 (n_1136, n1518);
  and g2014 (n1519, n847, n_1136);
  not g2015 (n_1137, n1519);
  and g2016 (n1520, n851, n_1137);
  not g2017 (n_1138, n1520);
  and g2018 (n1521, n855, n_1138);
  not g2019 (n_1139, n1521);
  and g2020 (n1522, n859, n_1139);
  not g2021 (n_1140, n1522);
  and g2022 (n1523, n863, n_1140);
  not g2023 (n_1141, n1523);
  and g2024 (n1524, n867, n_1141);
  not g2025 (n_1142, n1524);
  and g2026 (n1525, n871, n_1142);
  not g2027 (n_1143, n1525);
  and g2028 (n1526, n875, n_1143);
  not g2029 (n_1144, n1526);
  and g2030 (n1527, n879, n_1144);
  not g2031 (n_1145, n1527);
  and g2032 (n1528, n883, n_1145);
  not g2033 (n_1146, n1528);
  and g2034 (n1529, n887, n_1146);
  not g2035 (n_1147, n1529);
  and g2036 (n1530, n891, n_1147);
  not g2037 (n_1148, n1530);
  and g2038 (n1531, n895, n_1148);
  not g2039 (n_1149, n1531);
  and g2040 (n1532, n899, n_1149);
  not g2041 (n_1150, n1532);
  and g2042 (n1533, n903, n_1150);
  not g2043 (n_1151, n1533);
  and g2044 (n1534, n907, n_1151);
  not g2045 (n_1152, n1534);
  and g2046 (n1535, n911, n_1152);
  not g2047 (n_1153, n1535);
  and g2048 (n1536, n915, n_1153);
  not g2049 (n_1154, n1536);
  and g2050 (n1537, n919, n_1154);
  not g2051 (n_1155, n1537);
  and g2052 (n1538, n923, n_1155);
  not g2053 (n_1156, n1538);
  and g2054 (n1539, n927, n_1156);
  not g2055 (n_1157, n1539);
  and g2056 (n1540, n931, n_1157);
  not g2057 (n_1158, n1540);
  and g2058 (n1541, n935, n_1158);
  not g2059 (n_1159, n1541);
  and g2060 (n1542, n939, n_1159);
  not g2061 (n_1160, n1542);
  and g2062 (n1543, n943, n_1160);
  not g2063 (n_1161, n1543);
  and g2064 (n1544, n947, n_1161);
  not g2065 (n_1162, n1544);
  and g2066 (n1545, n951, n_1162);
  not g2067 (n_1163, n1545);
  and g2068 (n1546, n955, n_1163);
  not g2069 (n_1164, n1546);
  and g2070 (n1547, n959, n_1164);
  not g2071 (n_1165, n1547);
  and g2072 (n1548, n963, n_1165);
  not g2073 (n_1166, n1548);
  and g2074 (n1549, n967, n_1166);
  not g2075 (n_1167, n1549);
  and g2076 (n1550, n971, n_1167);
  not g2077 (n_1168, n1550);
  and g2078 (n1551, n975, n_1168);
  not g2079 (n_1169, n1551);
  and g2080 (n1552, n979, n_1169);
  not g2081 (n_1170, n1552);
  and g2082 (n1553, n983, n_1170);
  not g2083 (n_1171, n1553);
  and g2084 (n1554, n987, n_1171);
  not g2085 (n_1172, n1554);
  and g2086 (n1555, n991, n_1172);
  not g2087 (n_1173, n1555);
  and g2088 (n1556, n995, n_1173);
  not g2089 (n_1174, n1556);
  and g2090 (n1557, n999, n_1174);
  not g2091 (n_1175, n1557);
  and g2092 (n1558, n1003, n_1175);
  not g2093 (n_1176, n1558);
  and g2094 (n1559, n1007, n_1176);
  not g2095 (n_1177, n1559);
  and g2096 (n1560, n1011, n_1177);
  not g2097 (n_1178, n1560);
  and g2098 (n1561, n1015, n_1178);
  not g2099 (n_1179, n1561);
  and g2100 (n1562, n1019, n_1179);
  not g2101 (n_1180, n1562);
  and g2102 (n1563, n1023, n_1180);
  not g2103 (n_1181, n1563);
  and g2104 (n1564, n1027, n_1181);
  not g2105 (n_1182, n1564);
  and g2106 (n1565, n1031, n_1182);
  not g2107 (n_1183, n1565);
  and g2108 (n1566, n1035, n_1183);
  not g2109 (n_1184, n1566);
  and g2110 (n1567, n1039, n_1184);
  not g2111 (n_1185, n1567);
  and g2112 (n1568, n1043, n_1185);
  not g2113 (n_1186, n1568);
  and g2114 (n1569, n1047, n_1186);
  not g2115 (n_1187, n1569);
  and g2116 (n1570, n1051, n_1187);
  not g2117 (n_1188, n1570);
  and g2118 (n1571, n1055, n_1188);
  not g2119 (n_1189, n1571);
  and g2120 (n1572, n1059, n_1189);
  and g2121 (n1573, n_3, n_9);
  and g2122 (n1574, n_850, n1573);
  not g2123 (n_1190, n1572);
  and g2124 (n1575, n_1190, n1574);
  and g2125 (n1576, n_14, n726);
  not g2126 (n_1191, n1575);
  and g2127 (n1577, n_1191, n1576);
  and g2128 (n1578, n_14, \req[3] );
  not g2129 (n_1192, n1578);
  and g2130 (n1579, \req[4] , n_1192);
  not g2131 (n_1193, n1577);
  and g2132 (\grant[4] , n_1193, n1579);
  not g2133 (n_1194, n399);
  and g2134 (n1581, n_1194, n1071);
  not g2135 (n_1195, n1581);
  and g2136 (n1582, n1076, n_1195);
  not g2137 (n_1196, n1582);
  and g2138 (n1583, n1080, n_1196);
  not g2139 (n_1197, n1583);
  and g2140 (n1584, n1084, n_1197);
  not g2141 (n_1198, n1584);
  and g2142 (n1585, n1088, n_1198);
  not g2143 (n_1199, n1585);
  and g2144 (n1586, n1092, n_1199);
  not g2145 (n_1200, n1586);
  and g2146 (n1587, n1096, n_1200);
  not g2147 (n_1201, n1587);
  and g2148 (n1588, n1100, n_1201);
  not g2149 (n_1202, n1588);
  and g2150 (n1589, n1104, n_1202);
  not g2151 (n_1203, n1589);
  and g2152 (n1590, n1108, n_1203);
  not g2153 (n_1204, n1590);
  and g2154 (n1591, n1112, n_1204);
  not g2155 (n_1205, n1591);
  and g2156 (n1592, n1116, n_1205);
  not g2157 (n_1206, n1592);
  and g2158 (n1593, n1120, n_1206);
  not g2159 (n_1207, n1593);
  and g2160 (n1594, n1124, n_1207);
  not g2161 (n_1208, n1594);
  and g2162 (n1595, n1128, n_1208);
  not g2163 (n_1209, n1595);
  and g2164 (n1596, n1132, n_1209);
  not g2165 (n_1210, n1596);
  and g2166 (n1597, n1136, n_1210);
  not g2167 (n_1211, n1597);
  and g2168 (n1598, n1140, n_1211);
  not g2169 (n_1212, n1598);
  and g2170 (n1599, n1144, n_1212);
  not g2171 (n_1213, n1599);
  and g2172 (n1600, n1148, n_1213);
  not g2173 (n_1214, n1600);
  and g2174 (n1601, n1152, n_1214);
  not g2175 (n_1215, n1601);
  and g2176 (n1602, n1156, n_1215);
  not g2177 (n_1216, n1602);
  and g2178 (n1603, n1160, n_1216);
  not g2179 (n_1217, n1603);
  and g2180 (n1604, n1164, n_1217);
  not g2181 (n_1218, n1604);
  and g2182 (n1605, n1168, n_1218);
  not g2183 (n_1219, n1605);
  and g2184 (n1606, n1172, n_1219);
  not g2185 (n_1220, n1606);
  and g2186 (n1607, n1176, n_1220);
  not g2187 (n_1221, n1607);
  and g2188 (n1608, n1180, n_1221);
  not g2189 (n_1222, n1608);
  and g2190 (n1609, n1184, n_1222);
  not g2191 (n_1223, n1609);
  and g2192 (n1610, n1188, n_1223);
  not g2193 (n_1224, n1610);
  and g2194 (n1611, n1192, n_1224);
  not g2195 (n_1225, n1611);
  and g2196 (n1612, n1196, n_1225);
  not g2197 (n_1226, n1612);
  and g2198 (n1613, n1200, n_1226);
  not g2199 (n_1227, n1613);
  and g2200 (n1614, n1204, n_1227);
  not g2201 (n_1228, n1614);
  and g2202 (n1615, n1208, n_1228);
  not g2203 (n_1229, n1615);
  and g2204 (n1616, n1212, n_1229);
  not g2205 (n_1230, n1616);
  and g2206 (n1617, n1216, n_1230);
  not g2207 (n_1231, n1617);
  and g2208 (n1618, n1220, n_1231);
  not g2209 (n_1232, n1618);
  and g2210 (n1619, n1224, n_1232);
  not g2211 (n_1233, n1619);
  and g2212 (n1620, n1228, n_1233);
  not g2213 (n_1234, n1620);
  and g2214 (n1621, n1232, n_1234);
  not g2215 (n_1235, n1621);
  and g2216 (n1622, n1236, n_1235);
  not g2217 (n_1236, n1622);
  and g2218 (n1623, n1240, n_1236);
  not g2219 (n_1237, n1623);
  and g2220 (n1624, n1244, n_1237);
  not g2221 (n_1238, n1624);
  and g2222 (n1625, n1248, n_1238);
  not g2223 (n_1239, n1625);
  and g2224 (n1626, n1252, n_1239);
  not g2225 (n_1240, n1626);
  and g2226 (n1627, n1256, n_1240);
  not g2227 (n_1241, n1627);
  and g2228 (n1628, n1260, n_1241);
  not g2229 (n_1242, n1628);
  and g2230 (n1629, n1264, n_1242);
  not g2231 (n_1243, n1629);
  and g2232 (n1630, n1268, n_1243);
  not g2233 (n_1244, n1630);
  and g2234 (n1631, n1272, n_1244);
  not g2235 (n_1245, n1631);
  and g2236 (n1632, n1276, n_1245);
  not g2237 (n_1246, n1632);
  and g2238 (n1633, n1280, n_1246);
  not g2239 (n_1247, n1633);
  and g2240 (n1634, n1284, n_1247);
  not g2241 (n_1248, n1634);
  and g2242 (n1635, n1288, n_1248);
  not g2243 (n_1249, n1635);
  and g2244 (n1636, n1292, n_1249);
  not g2245 (n_1250, n1636);
  and g2246 (n1637, n1296, n_1250);
  not g2247 (n_1251, n1637);
  and g2248 (n1638, n1300, n_1251);
  not g2249 (n_1252, n1638);
  and g2250 (n1639, n1304, n_1252);
  not g2251 (n_1253, n1639);
  and g2252 (n1640, n1308, n_1253);
  not g2253 (n_1254, n1640);
  and g2254 (n1641, n1312, n_1254);
  not g2255 (n_1255, n1641);
  and g2256 (n1642, n1316, n_1255);
  not g2257 (n_1256, n1642);
  and g2258 (n1643, n1320, n_1256);
  not g2259 (n_1257, n1643);
  and g2260 (n1644, n1324, n_1257);
  not g2261 (n_1258, n1644);
  and g2262 (n1645, n1328, n_1258);
  not g2263 (n_1259, n1645);
  and g2264 (n1646, n1332, n_1259);
  not g2265 (n_1260, n1646);
  and g2266 (n1647, n1336, n_1260);
  not g2267 (n_1261, n1647);
  and g2268 (n1648, n1340, n_1261);
  not g2269 (n_1262, n1648);
  and g2270 (n1649, n1344, n_1262);
  not g2271 (n_1263, n1649);
  and g2272 (n1650, n1348, n_1263);
  not g2273 (n_1264, n1650);
  and g2274 (n1651, n1352, n_1264);
  not g2275 (n_1265, n1651);
  and g2276 (n1652, n1356, n_1265);
  not g2277 (n_1266, n1652);
  and g2278 (n1653, n1360, n_1266);
  not g2279 (n_1267, n1653);
  and g2280 (n1654, n1364, n_1267);
  not g2281 (n_1268, n1654);
  and g2282 (n1655, n1368, n_1268);
  not g2283 (n_1269, n1655);
  and g2284 (n1656, n1372, n_1269);
  not g2285 (n_1270, n1656);
  and g2286 (n1657, n1376, n_1270);
  not g2287 (n_1271, n1657);
  and g2288 (n1658, n1380, n_1271);
  not g2289 (n_1272, n1658);
  and g2290 (n1659, n1384, n_1272);
  not g2291 (n_1273, n1659);
  and g2292 (n1660, n1388, n_1273);
  not g2293 (n_1274, n1660);
  and g2294 (n1661, n1392, n_1274);
  not g2295 (n_1275, n1661);
  and g2296 (n1662, n1396, n_1275);
  and g2297 (n1663, n388, n_1020);
  not g2298 (n_1276, n1662);
  and g2299 (n1664, n_1276, n1663);
  not g2300 (n_1277, n1664);
  and g2301 (n1665, n392, n_1277);
  and g2302 (n1666, \req[5] , n_24);
  not g2303 (n_1278, n1665);
  and g2304 (\grant[5] , n_1278, n1666);
  not g2305 (n_1279, n738);
  and g2306 (n1668, n403, n_1279);
  not g2307 (n_1280, n1668);
  and g2308 (n1669, n408, n_1280);
  not g2309 (n_1281, n1669);
  and g2310 (n1670, n412, n_1281);
  not g2311 (n_1282, n1670);
  and g2312 (n1671, n416, n_1282);
  not g2313 (n_1283, n1671);
  and g2314 (n1672, n420, n_1283);
  not g2315 (n_1284, n1672);
  and g2316 (n1673, n424, n_1284);
  not g2317 (n_1285, n1673);
  and g2318 (n1674, n428, n_1285);
  not g2319 (n_1286, n1674);
  and g2320 (n1675, n432, n_1286);
  not g2321 (n_1287, n1675);
  and g2322 (n1676, n436, n_1287);
  not g2323 (n_1288, n1676);
  and g2324 (n1677, n440, n_1288);
  not g2325 (n_1289, n1677);
  and g2326 (n1678, n444, n_1289);
  not g2327 (n_1290, n1678);
  and g2328 (n1679, n448, n_1290);
  not g2329 (n_1291, n1679);
  and g2330 (n1680, n452, n_1291);
  not g2331 (n_1292, n1680);
  and g2332 (n1681, n456, n_1292);
  not g2333 (n_1293, n1681);
  and g2334 (n1682, n460, n_1293);
  not g2335 (n_1294, n1682);
  and g2336 (n1683, n464, n_1294);
  not g2337 (n_1295, n1683);
  and g2338 (n1684, n468, n_1295);
  not g2339 (n_1296, n1684);
  and g2340 (n1685, n472, n_1296);
  not g2341 (n_1297, n1685);
  and g2342 (n1686, n476, n_1297);
  not g2343 (n_1298, n1686);
  and g2344 (n1687, n480, n_1298);
  not g2345 (n_1299, n1687);
  and g2346 (n1688, n484, n_1299);
  not g2347 (n_1300, n1688);
  and g2348 (n1689, n488, n_1300);
  not g2349 (n_1301, n1689);
  and g2350 (n1690, n492, n_1301);
  not g2351 (n_1302, n1690);
  and g2352 (n1691, n496, n_1302);
  not g2353 (n_1303, n1691);
  and g2354 (n1692, n500, n_1303);
  not g2355 (n_1304, n1692);
  and g2356 (n1693, n504, n_1304);
  not g2357 (n_1305, n1693);
  and g2358 (n1694, n508, n_1305);
  not g2359 (n_1306, n1694);
  and g2360 (n1695, n512, n_1306);
  not g2361 (n_1307, n1695);
  and g2362 (n1696, n516, n_1307);
  not g2363 (n_1308, n1696);
  and g2364 (n1697, n520, n_1308);
  not g2365 (n_1309, n1697);
  and g2366 (n1698, n524, n_1309);
  not g2367 (n_1310, n1698);
  and g2368 (n1699, n528, n_1310);
  not g2369 (n_1311, n1699);
  and g2370 (n1700, n532, n_1311);
  not g2371 (n_1312, n1700);
  and g2372 (n1701, n536, n_1312);
  not g2373 (n_1313, n1701);
  and g2374 (n1702, n540, n_1313);
  not g2375 (n_1314, n1702);
  and g2376 (n1703, n544, n_1314);
  not g2377 (n_1315, n1703);
  and g2378 (n1704, n548, n_1315);
  not g2379 (n_1316, n1704);
  and g2380 (n1705, n552, n_1316);
  not g2381 (n_1317, n1705);
  and g2382 (n1706, n556, n_1317);
  not g2383 (n_1318, n1706);
  and g2384 (n1707, n560, n_1318);
  not g2385 (n_1319, n1707);
  and g2386 (n1708, n564, n_1319);
  not g2387 (n_1320, n1708);
  and g2388 (n1709, n568, n_1320);
  not g2389 (n_1321, n1709);
  and g2390 (n1710, n572, n_1321);
  not g2391 (n_1322, n1710);
  and g2392 (n1711, n576, n_1322);
  not g2393 (n_1323, n1711);
  and g2394 (n1712, n580, n_1323);
  not g2395 (n_1324, n1712);
  and g2396 (n1713, n584, n_1324);
  not g2397 (n_1325, n1713);
  and g2398 (n1714, n588, n_1325);
  not g2399 (n_1326, n1714);
  and g2400 (n1715, n592, n_1326);
  not g2401 (n_1327, n1715);
  and g2402 (n1716, n596, n_1327);
  not g2403 (n_1328, n1716);
  and g2404 (n1717, n600, n_1328);
  not g2405 (n_1329, n1717);
  and g2406 (n1718, n604, n_1329);
  not g2407 (n_1330, n1718);
  and g2408 (n1719, n608, n_1330);
  not g2409 (n_1331, n1719);
  and g2410 (n1720, n612, n_1331);
  not g2411 (n_1332, n1720);
  and g2412 (n1721, n616, n_1332);
  not g2413 (n_1333, n1721);
  and g2414 (n1722, n620, n_1333);
  not g2415 (n_1334, n1722);
  and g2416 (n1723, n624, n_1334);
  not g2417 (n_1335, n1723);
  and g2418 (n1724, n628, n_1335);
  not g2419 (n_1336, n1724);
  and g2420 (n1725, n632, n_1336);
  not g2421 (n_1337, n1725);
  and g2422 (n1726, n636, n_1337);
  not g2423 (n_1338, n1726);
  and g2424 (n1727, n640, n_1338);
  not g2425 (n_1339, n1727);
  and g2426 (n1728, n644, n_1339);
  not g2427 (n_1340, n1728);
  and g2428 (n1729, n648, n_1340);
  not g2429 (n_1341, n1729);
  and g2430 (n1730, n652, n_1341);
  not g2431 (n_1342, n1730);
  and g2432 (n1731, n656, n_1342);
  not g2433 (n_1343, n1731);
  and g2434 (n1732, n660, n_1343);
  not g2435 (n_1344, n1732);
  and g2436 (n1733, n664, n_1344);
  not g2437 (n_1345, n1733);
  and g2438 (n1734, n668, n_1345);
  not g2439 (n_1346, n1734);
  and g2440 (n1735, n672, n_1346);
  not g2441 (n_1347, n1735);
  and g2442 (n1736, n676, n_1347);
  not g2443 (n_1348, n1736);
  and g2444 (n1737, n680, n_1348);
  not g2445 (n_1349, n1737);
  and g2446 (n1738, n684, n_1349);
  not g2447 (n_1350, n1738);
  and g2448 (n1739, n688, n_1350);
  not g2449 (n_1351, n1739);
  and g2450 (n1740, n692, n_1351);
  not g2451 (n_1352, n1740);
  and g2452 (n1741, n696, n_1352);
  not g2453 (n_1353, n1741);
  and g2454 (n1742, n700, n_1353);
  not g2455 (n_1354, n1742);
  and g2456 (n1743, n704, n_1354);
  not g2457 (n_1355, n1743);
  and g2458 (n1744, n708, n_1355);
  not g2459 (n_1356, n1744);
  and g2460 (n1745, n712, n_1356);
  not g2461 (n_1357, n1745);
  and g2462 (n1746, n716, n_1357);
  not g2463 (n_1358, n1746);
  and g2464 (n1747, n720, n_1358);
  not g2465 (n_1359, n1747);
  and g2466 (n1748, n1484, n_1359);
  not g2467 (n_1360, n1748);
  and g2468 (n1749, n1486, n_1360);
  and g2469 (n1750, n727, n_1106);
  not g2470 (n_1361, n1749);
  and g2471 (n1751, n_1361, n1750);
  not g2472 (n_1362, n1751);
  and g2473 (n1752, n731, n_1362);
  and g2474 (n1753, \req[6] , n_605);
  not g2475 (n_1363, n1752);
  and g2476 (\grant[6] , n_1363, n1753);
  not g2477 (n_1364, n1075);
  and g2478 (n1755, n742, n_1364);
  not g2479 (n_1365, n1755);
  and g2480 (n1756, n747, n_1365);
  not g2481 (n_1366, n1756);
  and g2482 (n1757, n751, n_1366);
  not g2483 (n_1367, n1757);
  and g2484 (n1758, n755, n_1367);
  not g2485 (n_1368, n1758);
  and g2486 (n1759, n759, n_1368);
  not g2487 (n_1369, n1759);
  and g2488 (n1760, n763, n_1369);
  not g2489 (n_1370, n1760);
  and g2490 (n1761, n767, n_1370);
  not g2491 (n_1371, n1761);
  and g2492 (n1762, n771, n_1371);
  not g2493 (n_1372, n1762);
  and g2494 (n1763, n775, n_1372);
  not g2495 (n_1373, n1763);
  and g2496 (n1764, n779, n_1373);
  not g2497 (n_1374, n1764);
  and g2498 (n1765, n783, n_1374);
  not g2499 (n_1375, n1765);
  and g2500 (n1766, n787, n_1375);
  not g2501 (n_1376, n1766);
  and g2502 (n1767, n791, n_1376);
  not g2503 (n_1377, n1767);
  and g2504 (n1768, n795, n_1377);
  not g2505 (n_1378, n1768);
  and g2506 (n1769, n799, n_1378);
  not g2507 (n_1379, n1769);
  and g2508 (n1770, n803, n_1379);
  not g2509 (n_1380, n1770);
  and g2510 (n1771, n807, n_1380);
  not g2511 (n_1381, n1771);
  and g2512 (n1772, n811, n_1381);
  not g2513 (n_1382, n1772);
  and g2514 (n1773, n815, n_1382);
  not g2515 (n_1383, n1773);
  and g2516 (n1774, n819, n_1383);
  not g2517 (n_1384, n1774);
  and g2518 (n1775, n823, n_1384);
  not g2519 (n_1385, n1775);
  and g2520 (n1776, n827, n_1385);
  not g2521 (n_1386, n1776);
  and g2522 (n1777, n831, n_1386);
  not g2523 (n_1387, n1777);
  and g2524 (n1778, n835, n_1387);
  not g2525 (n_1388, n1778);
  and g2526 (n1779, n839, n_1388);
  not g2527 (n_1389, n1779);
  and g2528 (n1780, n843, n_1389);
  not g2529 (n_1390, n1780);
  and g2530 (n1781, n847, n_1390);
  not g2531 (n_1391, n1781);
  and g2532 (n1782, n851, n_1391);
  not g2533 (n_1392, n1782);
  and g2534 (n1783, n855, n_1392);
  not g2535 (n_1393, n1783);
  and g2536 (n1784, n859, n_1393);
  not g2537 (n_1394, n1784);
  and g2538 (n1785, n863, n_1394);
  not g2539 (n_1395, n1785);
  and g2540 (n1786, n867, n_1395);
  not g2541 (n_1396, n1786);
  and g2542 (n1787, n871, n_1396);
  not g2543 (n_1397, n1787);
  and g2544 (n1788, n875, n_1397);
  not g2545 (n_1398, n1788);
  and g2546 (n1789, n879, n_1398);
  not g2547 (n_1399, n1789);
  and g2548 (n1790, n883, n_1399);
  not g2549 (n_1400, n1790);
  and g2550 (n1791, n887, n_1400);
  not g2551 (n_1401, n1791);
  and g2552 (n1792, n891, n_1401);
  not g2553 (n_1402, n1792);
  and g2554 (n1793, n895, n_1402);
  not g2555 (n_1403, n1793);
  and g2556 (n1794, n899, n_1403);
  not g2557 (n_1404, n1794);
  and g2558 (n1795, n903, n_1404);
  not g2559 (n_1405, n1795);
  and g2560 (n1796, n907, n_1405);
  not g2561 (n_1406, n1796);
  and g2562 (n1797, n911, n_1406);
  not g2563 (n_1407, n1797);
  and g2564 (n1798, n915, n_1407);
  not g2565 (n_1408, n1798);
  and g2566 (n1799, n919, n_1408);
  not g2567 (n_1409, n1799);
  and g2568 (n1800, n923, n_1409);
  not g2569 (n_1410, n1800);
  and g2570 (n1801, n927, n_1410);
  not g2571 (n_1411, n1801);
  and g2572 (n1802, n931, n_1411);
  not g2573 (n_1412, n1802);
  and g2574 (n1803, n935, n_1412);
  not g2575 (n_1413, n1803);
  and g2576 (n1804, n939, n_1413);
  not g2577 (n_1414, n1804);
  and g2578 (n1805, n943, n_1414);
  not g2579 (n_1415, n1805);
  and g2580 (n1806, n947, n_1415);
  not g2581 (n_1416, n1806);
  and g2582 (n1807, n951, n_1416);
  not g2583 (n_1417, n1807);
  and g2584 (n1808, n955, n_1417);
  not g2585 (n_1418, n1808);
  and g2586 (n1809, n959, n_1418);
  not g2587 (n_1419, n1809);
  and g2588 (n1810, n963, n_1419);
  not g2589 (n_1420, n1810);
  and g2590 (n1811, n967, n_1420);
  not g2591 (n_1421, n1811);
  and g2592 (n1812, n971, n_1421);
  not g2593 (n_1422, n1812);
  and g2594 (n1813, n975, n_1422);
  not g2595 (n_1423, n1813);
  and g2596 (n1814, n979, n_1423);
  not g2597 (n_1424, n1814);
  and g2598 (n1815, n983, n_1424);
  not g2599 (n_1425, n1815);
  and g2600 (n1816, n987, n_1425);
  not g2601 (n_1426, n1816);
  and g2602 (n1817, n991, n_1426);
  not g2603 (n_1427, n1817);
  and g2604 (n1818, n995, n_1427);
  not g2605 (n_1428, n1818);
  and g2606 (n1819, n999, n_1428);
  not g2607 (n_1429, n1819);
  and g2608 (n1820, n1003, n_1429);
  not g2609 (n_1430, n1820);
  and g2610 (n1821, n1007, n_1430);
  not g2611 (n_1431, n1821);
  and g2612 (n1822, n1011, n_1431);
  not g2613 (n_1432, n1822);
  and g2614 (n1823, n1015, n_1432);
  not g2615 (n_1433, n1823);
  and g2616 (n1824, n1019, n_1433);
  not g2617 (n_1434, n1824);
  and g2618 (n1825, n1023, n_1434);
  not g2619 (n_1435, n1825);
  and g2620 (n1826, n1027, n_1435);
  not g2621 (n_1436, n1826);
  and g2622 (n1827, n1031, n_1436);
  not g2623 (n_1437, n1827);
  and g2624 (n1828, n1035, n_1437);
  not g2625 (n_1438, n1828);
  and g2626 (n1829, n1039, n_1438);
  not g2627 (n_1439, n1829);
  and g2628 (n1830, n1043, n_1439);
  not g2629 (n_1440, n1830);
  and g2630 (n1831, n1047, n_1440);
  not g2631 (n_1441, n1831);
  and g2632 (n1832, n1051, n_1441);
  not g2633 (n_1442, n1832);
  and g2634 (n1833, n1055, n_1442);
  not g2635 (n_1443, n1833);
  and g2636 (n1834, n1059, n_1443);
  not g2637 (n_1444, n1834);
  and g2638 (n1835, n1574, n_1444);
  not g2639 (n_1445, n1835);
  and g2640 (n1836, n1576, n_1445);
  and g2641 (n1837, n1064, n_1192);
  not g2642 (n_1446, n1836);
  and g2643 (n1838, n_1446, n1837);
  not g2644 (n_1447, n1838);
  and g2645 (n1839, n1068, n_1447);
  and g2646 (n1840, \req[7] , n_855);
  not g2647 (n_1448, n1839);
  and g2648 (\grant[7] , n_1448, n1840);
  not g2649 (n_1449, n407);
  and g2650 (n1842, n_1449, n1079);
  not g2651 (n_1450, n1842);
  and g2652 (n1843, n1084, n_1450);
  not g2653 (n_1451, n1843);
  and g2654 (n1844, n1088, n_1451);
  not g2655 (n_1452, n1844);
  and g2656 (n1845, n1092, n_1452);
  not g2657 (n_1453, n1845);
  and g2658 (n1846, n1096, n_1453);
  not g2659 (n_1454, n1846);
  and g2660 (n1847, n1100, n_1454);
  not g2661 (n_1455, n1847);
  and g2662 (n1848, n1104, n_1455);
  not g2663 (n_1456, n1848);
  and g2664 (n1849, n1108, n_1456);
  not g2665 (n_1457, n1849);
  and g2666 (n1850, n1112, n_1457);
  not g2667 (n_1458, n1850);
  and g2668 (n1851, n1116, n_1458);
  not g2669 (n_1459, n1851);
  and g2670 (n1852, n1120, n_1459);
  not g2671 (n_1460, n1852);
  and g2672 (n1853, n1124, n_1460);
  not g2673 (n_1461, n1853);
  and g2674 (n1854, n1128, n_1461);
  not g2675 (n_1462, n1854);
  and g2676 (n1855, n1132, n_1462);
  not g2677 (n_1463, n1855);
  and g2678 (n1856, n1136, n_1463);
  not g2679 (n_1464, n1856);
  and g2680 (n1857, n1140, n_1464);
  not g2681 (n_1465, n1857);
  and g2682 (n1858, n1144, n_1465);
  not g2683 (n_1466, n1858);
  and g2684 (n1859, n1148, n_1466);
  not g2685 (n_1467, n1859);
  and g2686 (n1860, n1152, n_1467);
  not g2687 (n_1468, n1860);
  and g2688 (n1861, n1156, n_1468);
  not g2689 (n_1469, n1861);
  and g2690 (n1862, n1160, n_1469);
  not g2691 (n_1470, n1862);
  and g2692 (n1863, n1164, n_1470);
  not g2693 (n_1471, n1863);
  and g2694 (n1864, n1168, n_1471);
  not g2695 (n_1472, n1864);
  and g2696 (n1865, n1172, n_1472);
  not g2697 (n_1473, n1865);
  and g2698 (n1866, n1176, n_1473);
  not g2699 (n_1474, n1866);
  and g2700 (n1867, n1180, n_1474);
  not g2701 (n_1475, n1867);
  and g2702 (n1868, n1184, n_1475);
  not g2703 (n_1476, n1868);
  and g2704 (n1869, n1188, n_1476);
  not g2705 (n_1477, n1869);
  and g2706 (n1870, n1192, n_1477);
  not g2707 (n_1478, n1870);
  and g2708 (n1871, n1196, n_1478);
  not g2709 (n_1479, n1871);
  and g2710 (n1872, n1200, n_1479);
  not g2711 (n_1480, n1872);
  and g2712 (n1873, n1204, n_1480);
  not g2713 (n_1481, n1873);
  and g2714 (n1874, n1208, n_1481);
  not g2715 (n_1482, n1874);
  and g2716 (n1875, n1212, n_1482);
  not g2717 (n_1483, n1875);
  and g2718 (n1876, n1216, n_1483);
  not g2719 (n_1484, n1876);
  and g2720 (n1877, n1220, n_1484);
  not g2721 (n_1485, n1877);
  and g2722 (n1878, n1224, n_1485);
  not g2723 (n_1486, n1878);
  and g2724 (n1879, n1228, n_1486);
  not g2725 (n_1487, n1879);
  and g2726 (n1880, n1232, n_1487);
  not g2727 (n_1488, n1880);
  and g2728 (n1881, n1236, n_1488);
  not g2729 (n_1489, n1881);
  and g2730 (n1882, n1240, n_1489);
  not g2731 (n_1490, n1882);
  and g2732 (n1883, n1244, n_1490);
  not g2733 (n_1491, n1883);
  and g2734 (n1884, n1248, n_1491);
  not g2735 (n_1492, n1884);
  and g2736 (n1885, n1252, n_1492);
  not g2737 (n_1493, n1885);
  and g2738 (n1886, n1256, n_1493);
  not g2739 (n_1494, n1886);
  and g2740 (n1887, n1260, n_1494);
  not g2741 (n_1495, n1887);
  and g2742 (n1888, n1264, n_1495);
  not g2743 (n_1496, n1888);
  and g2744 (n1889, n1268, n_1496);
  not g2745 (n_1497, n1889);
  and g2746 (n1890, n1272, n_1497);
  not g2747 (n_1498, n1890);
  and g2748 (n1891, n1276, n_1498);
  not g2749 (n_1499, n1891);
  and g2750 (n1892, n1280, n_1499);
  not g2751 (n_1500, n1892);
  and g2752 (n1893, n1284, n_1500);
  not g2753 (n_1501, n1893);
  and g2754 (n1894, n1288, n_1501);
  not g2755 (n_1502, n1894);
  and g2756 (n1895, n1292, n_1502);
  not g2757 (n_1503, n1895);
  and g2758 (n1896, n1296, n_1503);
  not g2759 (n_1504, n1896);
  and g2760 (n1897, n1300, n_1504);
  not g2761 (n_1505, n1897);
  and g2762 (n1898, n1304, n_1505);
  not g2763 (n_1506, n1898);
  and g2764 (n1899, n1308, n_1506);
  not g2765 (n_1507, n1899);
  and g2766 (n1900, n1312, n_1507);
  not g2767 (n_1508, n1900);
  and g2768 (n1901, n1316, n_1508);
  not g2769 (n_1509, n1901);
  and g2770 (n1902, n1320, n_1509);
  not g2771 (n_1510, n1902);
  and g2772 (n1903, n1324, n_1510);
  not g2773 (n_1511, n1903);
  and g2774 (n1904, n1328, n_1511);
  not g2775 (n_1512, n1904);
  and g2776 (n1905, n1332, n_1512);
  not g2777 (n_1513, n1905);
  and g2778 (n1906, n1336, n_1513);
  not g2779 (n_1514, n1906);
  and g2780 (n1907, n1340, n_1514);
  not g2781 (n_1515, n1907);
  and g2782 (n1908, n1344, n_1515);
  not g2783 (n_1516, n1908);
  and g2784 (n1909, n1348, n_1516);
  not g2785 (n_1517, n1909);
  and g2786 (n1910, n1352, n_1517);
  not g2787 (n_1518, n1910);
  and g2788 (n1911, n1356, n_1518);
  not g2789 (n_1519, n1911);
  and g2790 (n1912, n1360, n_1519);
  not g2791 (n_1520, n1912);
  and g2792 (n1913, n1364, n_1520);
  not g2793 (n_1521, n1913);
  and g2794 (n1914, n1368, n_1521);
  not g2795 (n_1522, n1914);
  and g2796 (n1915, n1372, n_1522);
  not g2797 (n_1523, n1915);
  and g2798 (n1916, n1376, n_1523);
  not g2799 (n_1524, n1916);
  and g2800 (n1917, n1380, n_1524);
  not g2801 (n_1525, n1917);
  and g2802 (n1918, n1384, n_1525);
  not g2803 (n_1526, n1918);
  and g2804 (n1919, n1388, n_1526);
  not g2805 (n_1527, n1919);
  and g2806 (n1920, n1392, n_1527);
  not g2807 (n_1528, n1920);
  and g2808 (n1921, n1396, n_1528);
  not g2809 (n_1529, n1921);
  and g2810 (n1922, n1663, n_1529);
  not g2811 (n_1530, n1922);
  and g2812 (n1923, n392, n_1530);
  not g2813 (n_1531, n1923);
  and g2814 (n1924, n396, n_1531);
  not g2815 (n_1532, n1924);
  and g2816 (n1925, n400, n_1532);
  and g2817 (n1926, \req[8] , n_38);
  not g2818 (n_1533, n1925);
  and g2819 (\grant[8] , n_1533, n1926);
  not g2820 (n_1534, n746);
  and g2821 (n1928, n411, n_1534);
  not g2822 (n_1535, n1928);
  and g2823 (n1929, n416, n_1535);
  not g2824 (n_1536, n1929);
  and g2825 (n1930, n420, n_1536);
  not g2826 (n_1537, n1930);
  and g2827 (n1931, n424, n_1537);
  not g2828 (n_1538, n1931);
  and g2829 (n1932, n428, n_1538);
  not g2830 (n_1539, n1932);
  and g2831 (n1933, n432, n_1539);
  not g2832 (n_1540, n1933);
  and g2833 (n1934, n436, n_1540);
  not g2834 (n_1541, n1934);
  and g2835 (n1935, n440, n_1541);
  not g2836 (n_1542, n1935);
  and g2837 (n1936, n444, n_1542);
  not g2838 (n_1543, n1936);
  and g2839 (n1937, n448, n_1543);
  not g2840 (n_1544, n1937);
  and g2841 (n1938, n452, n_1544);
  not g2842 (n_1545, n1938);
  and g2843 (n1939, n456, n_1545);
  not g2844 (n_1546, n1939);
  and g2845 (n1940, n460, n_1546);
  not g2846 (n_1547, n1940);
  and g2847 (n1941, n464, n_1547);
  not g2848 (n_1548, n1941);
  and g2849 (n1942, n468, n_1548);
  not g2850 (n_1549, n1942);
  and g2851 (n1943, n472, n_1549);
  not g2852 (n_1550, n1943);
  and g2853 (n1944, n476, n_1550);
  not g2854 (n_1551, n1944);
  and g2855 (n1945, n480, n_1551);
  not g2856 (n_1552, n1945);
  and g2857 (n1946, n484, n_1552);
  not g2858 (n_1553, n1946);
  and g2859 (n1947, n488, n_1553);
  not g2860 (n_1554, n1947);
  and g2861 (n1948, n492, n_1554);
  not g2862 (n_1555, n1948);
  and g2863 (n1949, n496, n_1555);
  not g2864 (n_1556, n1949);
  and g2865 (n1950, n500, n_1556);
  not g2866 (n_1557, n1950);
  and g2867 (n1951, n504, n_1557);
  not g2868 (n_1558, n1951);
  and g2869 (n1952, n508, n_1558);
  not g2870 (n_1559, n1952);
  and g2871 (n1953, n512, n_1559);
  not g2872 (n_1560, n1953);
  and g2873 (n1954, n516, n_1560);
  not g2874 (n_1561, n1954);
  and g2875 (n1955, n520, n_1561);
  not g2876 (n_1562, n1955);
  and g2877 (n1956, n524, n_1562);
  not g2878 (n_1563, n1956);
  and g2879 (n1957, n528, n_1563);
  not g2880 (n_1564, n1957);
  and g2881 (n1958, n532, n_1564);
  not g2882 (n_1565, n1958);
  and g2883 (n1959, n536, n_1565);
  not g2884 (n_1566, n1959);
  and g2885 (n1960, n540, n_1566);
  not g2886 (n_1567, n1960);
  and g2887 (n1961, n544, n_1567);
  not g2888 (n_1568, n1961);
  and g2889 (n1962, n548, n_1568);
  not g2890 (n_1569, n1962);
  and g2891 (n1963, n552, n_1569);
  not g2892 (n_1570, n1963);
  and g2893 (n1964, n556, n_1570);
  not g2894 (n_1571, n1964);
  and g2895 (n1965, n560, n_1571);
  not g2896 (n_1572, n1965);
  and g2897 (n1966, n564, n_1572);
  not g2898 (n_1573, n1966);
  and g2899 (n1967, n568, n_1573);
  not g2900 (n_1574, n1967);
  and g2901 (n1968, n572, n_1574);
  not g2902 (n_1575, n1968);
  and g2903 (n1969, n576, n_1575);
  not g2904 (n_1576, n1969);
  and g2905 (n1970, n580, n_1576);
  not g2906 (n_1577, n1970);
  and g2907 (n1971, n584, n_1577);
  not g2908 (n_1578, n1971);
  and g2909 (n1972, n588, n_1578);
  not g2910 (n_1579, n1972);
  and g2911 (n1973, n592, n_1579);
  not g2912 (n_1580, n1973);
  and g2913 (n1974, n596, n_1580);
  not g2914 (n_1581, n1974);
  and g2915 (n1975, n600, n_1581);
  not g2916 (n_1582, n1975);
  and g2917 (n1976, n604, n_1582);
  not g2918 (n_1583, n1976);
  and g2919 (n1977, n608, n_1583);
  not g2920 (n_1584, n1977);
  and g2921 (n1978, n612, n_1584);
  not g2922 (n_1585, n1978);
  and g2923 (n1979, n616, n_1585);
  not g2924 (n_1586, n1979);
  and g2925 (n1980, n620, n_1586);
  not g2926 (n_1587, n1980);
  and g2927 (n1981, n624, n_1587);
  not g2928 (n_1588, n1981);
  and g2929 (n1982, n628, n_1588);
  not g2930 (n_1589, n1982);
  and g2931 (n1983, n632, n_1589);
  not g2932 (n_1590, n1983);
  and g2933 (n1984, n636, n_1590);
  not g2934 (n_1591, n1984);
  and g2935 (n1985, n640, n_1591);
  not g2936 (n_1592, n1985);
  and g2937 (n1986, n644, n_1592);
  not g2938 (n_1593, n1986);
  and g2939 (n1987, n648, n_1593);
  not g2940 (n_1594, n1987);
  and g2941 (n1988, n652, n_1594);
  not g2942 (n_1595, n1988);
  and g2943 (n1989, n656, n_1595);
  not g2944 (n_1596, n1989);
  and g2945 (n1990, n660, n_1596);
  not g2946 (n_1597, n1990);
  and g2947 (n1991, n664, n_1597);
  not g2948 (n_1598, n1991);
  and g2949 (n1992, n668, n_1598);
  not g2950 (n_1599, n1992);
  and g2951 (n1993, n672, n_1599);
  not g2952 (n_1600, n1993);
  and g2953 (n1994, n676, n_1600);
  not g2954 (n_1601, n1994);
  and g2955 (n1995, n680, n_1601);
  not g2956 (n_1602, n1995);
  and g2957 (n1996, n684, n_1602);
  not g2958 (n_1603, n1996);
  and g2959 (n1997, n688, n_1603);
  not g2960 (n_1604, n1997);
  and g2961 (n1998, n692, n_1604);
  not g2962 (n_1605, n1998);
  and g2963 (n1999, n696, n_1605);
  not g2964 (n_1606, n1999);
  and g2965 (n2000, n700, n_1606);
  not g2966 (n_1607, n2000);
  and g2967 (n2001, n704, n_1607);
  not g2968 (n_1608, n2001);
  and g2969 (n2002, n708, n_1608);
  not g2970 (n_1609, n2002);
  and g2971 (n2003, n712, n_1609);
  not g2972 (n_1610, n2003);
  and g2973 (n2004, n716, n_1610);
  not g2974 (n_1611, n2004);
  and g2975 (n2005, n720, n_1611);
  not g2976 (n_1612, n2005);
  and g2977 (n2006, n1484, n_1612);
  not g2978 (n_1613, n2006);
  and g2979 (n2007, n1486, n_1613);
  not g2980 (n_1614, n2007);
  and g2981 (n2008, n1750, n_1614);
  not g2982 (n_1615, n2008);
  and g2983 (n2009, n731, n_1615);
  not g2984 (n_1616, n2009);
  and g2985 (n2010, n735, n_1616);
  not g2986 (n_1617, n2010);
  and g2987 (n2011, n739, n_1617);
  and g2988 (n2012, \req[9] , n_611);
  not g2989 (n_1618, n2011);
  and g2990 (\grant[9] , n_1618, n2012);
  not g2991 (n_1619, n1083);
  and g2992 (n2014, n750, n_1619);
  not g2993 (n_1620, n2014);
  and g2994 (n2015, n755, n_1620);
  not g2995 (n_1621, n2015);
  and g2996 (n2016, n759, n_1621);
  not g2997 (n_1622, n2016);
  and g2998 (n2017, n763, n_1622);
  not g2999 (n_1623, n2017);
  and g3000 (n2018, n767, n_1623);
  not g3001 (n_1624, n2018);
  and g3002 (n2019, n771, n_1624);
  not g3003 (n_1625, n2019);
  and g3004 (n2020, n775, n_1625);
  not g3005 (n_1626, n2020);
  and g3006 (n2021, n779, n_1626);
  not g3007 (n_1627, n2021);
  and g3008 (n2022, n783, n_1627);
  not g3009 (n_1628, n2022);
  and g3010 (n2023, n787, n_1628);
  not g3011 (n_1629, n2023);
  and g3012 (n2024, n791, n_1629);
  not g3013 (n_1630, n2024);
  and g3014 (n2025, n795, n_1630);
  not g3015 (n_1631, n2025);
  and g3016 (n2026, n799, n_1631);
  not g3017 (n_1632, n2026);
  and g3018 (n2027, n803, n_1632);
  not g3019 (n_1633, n2027);
  and g3020 (n2028, n807, n_1633);
  not g3021 (n_1634, n2028);
  and g3022 (n2029, n811, n_1634);
  not g3023 (n_1635, n2029);
  and g3024 (n2030, n815, n_1635);
  not g3025 (n_1636, n2030);
  and g3026 (n2031, n819, n_1636);
  not g3027 (n_1637, n2031);
  and g3028 (n2032, n823, n_1637);
  not g3029 (n_1638, n2032);
  and g3030 (n2033, n827, n_1638);
  not g3031 (n_1639, n2033);
  and g3032 (n2034, n831, n_1639);
  not g3033 (n_1640, n2034);
  and g3034 (n2035, n835, n_1640);
  not g3035 (n_1641, n2035);
  and g3036 (n2036, n839, n_1641);
  not g3037 (n_1642, n2036);
  and g3038 (n2037, n843, n_1642);
  not g3039 (n_1643, n2037);
  and g3040 (n2038, n847, n_1643);
  not g3041 (n_1644, n2038);
  and g3042 (n2039, n851, n_1644);
  not g3043 (n_1645, n2039);
  and g3044 (n2040, n855, n_1645);
  not g3045 (n_1646, n2040);
  and g3046 (n2041, n859, n_1646);
  not g3047 (n_1647, n2041);
  and g3048 (n2042, n863, n_1647);
  not g3049 (n_1648, n2042);
  and g3050 (n2043, n867, n_1648);
  not g3051 (n_1649, n2043);
  and g3052 (n2044, n871, n_1649);
  not g3053 (n_1650, n2044);
  and g3054 (n2045, n875, n_1650);
  not g3055 (n_1651, n2045);
  and g3056 (n2046, n879, n_1651);
  not g3057 (n_1652, n2046);
  and g3058 (n2047, n883, n_1652);
  not g3059 (n_1653, n2047);
  and g3060 (n2048, n887, n_1653);
  not g3061 (n_1654, n2048);
  and g3062 (n2049, n891, n_1654);
  not g3063 (n_1655, n2049);
  and g3064 (n2050, n895, n_1655);
  not g3065 (n_1656, n2050);
  and g3066 (n2051, n899, n_1656);
  not g3067 (n_1657, n2051);
  and g3068 (n2052, n903, n_1657);
  not g3069 (n_1658, n2052);
  and g3070 (n2053, n907, n_1658);
  not g3071 (n_1659, n2053);
  and g3072 (n2054, n911, n_1659);
  not g3073 (n_1660, n2054);
  and g3074 (n2055, n915, n_1660);
  not g3075 (n_1661, n2055);
  and g3076 (n2056, n919, n_1661);
  not g3077 (n_1662, n2056);
  and g3078 (n2057, n923, n_1662);
  not g3079 (n_1663, n2057);
  and g3080 (n2058, n927, n_1663);
  not g3081 (n_1664, n2058);
  and g3082 (n2059, n931, n_1664);
  not g3083 (n_1665, n2059);
  and g3084 (n2060, n935, n_1665);
  not g3085 (n_1666, n2060);
  and g3086 (n2061, n939, n_1666);
  not g3087 (n_1667, n2061);
  and g3088 (n2062, n943, n_1667);
  not g3089 (n_1668, n2062);
  and g3090 (n2063, n947, n_1668);
  not g3091 (n_1669, n2063);
  and g3092 (n2064, n951, n_1669);
  not g3093 (n_1670, n2064);
  and g3094 (n2065, n955, n_1670);
  not g3095 (n_1671, n2065);
  and g3096 (n2066, n959, n_1671);
  not g3097 (n_1672, n2066);
  and g3098 (n2067, n963, n_1672);
  not g3099 (n_1673, n2067);
  and g3100 (n2068, n967, n_1673);
  not g3101 (n_1674, n2068);
  and g3102 (n2069, n971, n_1674);
  not g3103 (n_1675, n2069);
  and g3104 (n2070, n975, n_1675);
  not g3105 (n_1676, n2070);
  and g3106 (n2071, n979, n_1676);
  not g3107 (n_1677, n2071);
  and g3108 (n2072, n983, n_1677);
  not g3109 (n_1678, n2072);
  and g3110 (n2073, n987, n_1678);
  not g3111 (n_1679, n2073);
  and g3112 (n2074, n991, n_1679);
  not g3113 (n_1680, n2074);
  and g3114 (n2075, n995, n_1680);
  not g3115 (n_1681, n2075);
  and g3116 (n2076, n999, n_1681);
  not g3117 (n_1682, n2076);
  and g3118 (n2077, n1003, n_1682);
  not g3119 (n_1683, n2077);
  and g3120 (n2078, n1007, n_1683);
  not g3121 (n_1684, n2078);
  and g3122 (n2079, n1011, n_1684);
  not g3123 (n_1685, n2079);
  and g3124 (n2080, n1015, n_1685);
  not g3125 (n_1686, n2080);
  and g3126 (n2081, n1019, n_1686);
  not g3127 (n_1687, n2081);
  and g3128 (n2082, n1023, n_1687);
  not g3129 (n_1688, n2082);
  and g3130 (n2083, n1027, n_1688);
  not g3131 (n_1689, n2083);
  and g3132 (n2084, n1031, n_1689);
  not g3133 (n_1690, n2084);
  and g3134 (n2085, n1035, n_1690);
  not g3135 (n_1691, n2085);
  and g3136 (n2086, n1039, n_1691);
  not g3137 (n_1692, n2086);
  and g3138 (n2087, n1043, n_1692);
  not g3139 (n_1693, n2087);
  and g3140 (n2088, n1047, n_1693);
  not g3141 (n_1694, n2088);
  and g3142 (n2089, n1051, n_1694);
  not g3143 (n_1695, n2089);
  and g3144 (n2090, n1055, n_1695);
  not g3145 (n_1696, n2090);
  and g3146 (n2091, n1059, n_1696);
  not g3147 (n_1697, n2091);
  and g3148 (n2092, n1574, n_1697);
  not g3149 (n_1698, n2092);
  and g3150 (n2093, n1576, n_1698);
  not g3151 (n_1699, n2093);
  and g3152 (n2094, n1837, n_1699);
  not g3153 (n_1700, n2094);
  and g3154 (n2095, n1068, n_1700);
  not g3155 (n_1701, n2095);
  and g3156 (n2096, n1072, n_1701);
  not g3157 (n_1702, n2096);
  and g3158 (n2097, n1076, n_1702);
  and g3159 (n2098, \req[10] , n_859);
  not g3160 (n_1703, n2097);
  and g3161 (\grant[10] , n_1703, n2098);
  not g3162 (n_1704, n415);
  and g3163 (n2100, n_1704, n1087);
  not g3164 (n_1705, n2100);
  and g3165 (n2101, n1092, n_1705);
  not g3166 (n_1706, n2101);
  and g3167 (n2102, n1096, n_1706);
  not g3168 (n_1707, n2102);
  and g3169 (n2103, n1100, n_1707);
  not g3170 (n_1708, n2103);
  and g3171 (n2104, n1104, n_1708);
  not g3172 (n_1709, n2104);
  and g3173 (n2105, n1108, n_1709);
  not g3174 (n_1710, n2105);
  and g3175 (n2106, n1112, n_1710);
  not g3176 (n_1711, n2106);
  and g3177 (n2107, n1116, n_1711);
  not g3178 (n_1712, n2107);
  and g3179 (n2108, n1120, n_1712);
  not g3180 (n_1713, n2108);
  and g3181 (n2109, n1124, n_1713);
  not g3182 (n_1714, n2109);
  and g3183 (n2110, n1128, n_1714);
  not g3184 (n_1715, n2110);
  and g3185 (n2111, n1132, n_1715);
  not g3186 (n_1716, n2111);
  and g3187 (n2112, n1136, n_1716);
  not g3188 (n_1717, n2112);
  and g3189 (n2113, n1140, n_1717);
  not g3190 (n_1718, n2113);
  and g3191 (n2114, n1144, n_1718);
  not g3192 (n_1719, n2114);
  and g3193 (n2115, n1148, n_1719);
  not g3194 (n_1720, n2115);
  and g3195 (n2116, n1152, n_1720);
  not g3196 (n_1721, n2116);
  and g3197 (n2117, n1156, n_1721);
  not g3198 (n_1722, n2117);
  and g3199 (n2118, n1160, n_1722);
  not g3200 (n_1723, n2118);
  and g3201 (n2119, n1164, n_1723);
  not g3202 (n_1724, n2119);
  and g3203 (n2120, n1168, n_1724);
  not g3204 (n_1725, n2120);
  and g3205 (n2121, n1172, n_1725);
  not g3206 (n_1726, n2121);
  and g3207 (n2122, n1176, n_1726);
  not g3208 (n_1727, n2122);
  and g3209 (n2123, n1180, n_1727);
  not g3210 (n_1728, n2123);
  and g3211 (n2124, n1184, n_1728);
  not g3212 (n_1729, n2124);
  and g3213 (n2125, n1188, n_1729);
  not g3214 (n_1730, n2125);
  and g3215 (n2126, n1192, n_1730);
  not g3216 (n_1731, n2126);
  and g3217 (n2127, n1196, n_1731);
  not g3218 (n_1732, n2127);
  and g3219 (n2128, n1200, n_1732);
  not g3220 (n_1733, n2128);
  and g3221 (n2129, n1204, n_1733);
  not g3222 (n_1734, n2129);
  and g3223 (n2130, n1208, n_1734);
  not g3224 (n_1735, n2130);
  and g3225 (n2131, n1212, n_1735);
  not g3226 (n_1736, n2131);
  and g3227 (n2132, n1216, n_1736);
  not g3228 (n_1737, n2132);
  and g3229 (n2133, n1220, n_1737);
  not g3230 (n_1738, n2133);
  and g3231 (n2134, n1224, n_1738);
  not g3232 (n_1739, n2134);
  and g3233 (n2135, n1228, n_1739);
  not g3234 (n_1740, n2135);
  and g3235 (n2136, n1232, n_1740);
  not g3236 (n_1741, n2136);
  and g3237 (n2137, n1236, n_1741);
  not g3238 (n_1742, n2137);
  and g3239 (n2138, n1240, n_1742);
  not g3240 (n_1743, n2138);
  and g3241 (n2139, n1244, n_1743);
  not g3242 (n_1744, n2139);
  and g3243 (n2140, n1248, n_1744);
  not g3244 (n_1745, n2140);
  and g3245 (n2141, n1252, n_1745);
  not g3246 (n_1746, n2141);
  and g3247 (n2142, n1256, n_1746);
  not g3248 (n_1747, n2142);
  and g3249 (n2143, n1260, n_1747);
  not g3250 (n_1748, n2143);
  and g3251 (n2144, n1264, n_1748);
  not g3252 (n_1749, n2144);
  and g3253 (n2145, n1268, n_1749);
  not g3254 (n_1750, n2145);
  and g3255 (n2146, n1272, n_1750);
  not g3256 (n_1751, n2146);
  and g3257 (n2147, n1276, n_1751);
  not g3258 (n_1752, n2147);
  and g3259 (n2148, n1280, n_1752);
  not g3260 (n_1753, n2148);
  and g3261 (n2149, n1284, n_1753);
  not g3262 (n_1754, n2149);
  and g3263 (n2150, n1288, n_1754);
  not g3264 (n_1755, n2150);
  and g3265 (n2151, n1292, n_1755);
  not g3266 (n_1756, n2151);
  and g3267 (n2152, n1296, n_1756);
  not g3268 (n_1757, n2152);
  and g3269 (n2153, n1300, n_1757);
  not g3270 (n_1758, n2153);
  and g3271 (n2154, n1304, n_1758);
  not g3272 (n_1759, n2154);
  and g3273 (n2155, n1308, n_1759);
  not g3274 (n_1760, n2155);
  and g3275 (n2156, n1312, n_1760);
  not g3276 (n_1761, n2156);
  and g3277 (n2157, n1316, n_1761);
  not g3278 (n_1762, n2157);
  and g3279 (n2158, n1320, n_1762);
  not g3280 (n_1763, n2158);
  and g3281 (n2159, n1324, n_1763);
  not g3282 (n_1764, n2159);
  and g3283 (n2160, n1328, n_1764);
  not g3284 (n_1765, n2160);
  and g3285 (n2161, n1332, n_1765);
  not g3286 (n_1766, n2161);
  and g3287 (n2162, n1336, n_1766);
  not g3288 (n_1767, n2162);
  and g3289 (n2163, n1340, n_1767);
  not g3290 (n_1768, n2163);
  and g3291 (n2164, n1344, n_1768);
  not g3292 (n_1769, n2164);
  and g3293 (n2165, n1348, n_1769);
  not g3294 (n_1770, n2165);
  and g3295 (n2166, n1352, n_1770);
  not g3296 (n_1771, n2166);
  and g3297 (n2167, n1356, n_1771);
  not g3298 (n_1772, n2167);
  and g3299 (n2168, n1360, n_1772);
  not g3300 (n_1773, n2168);
  and g3301 (n2169, n1364, n_1773);
  not g3302 (n_1774, n2169);
  and g3303 (n2170, n1368, n_1774);
  not g3304 (n_1775, n2170);
  and g3305 (n2171, n1372, n_1775);
  not g3306 (n_1776, n2171);
  and g3307 (n2172, n1376, n_1776);
  not g3308 (n_1777, n2172);
  and g3309 (n2173, n1380, n_1777);
  not g3310 (n_1778, n2173);
  and g3311 (n2174, n1384, n_1778);
  not g3312 (n_1779, n2174);
  and g3313 (n2175, n1388, n_1779);
  not g3314 (n_1780, n2175);
  and g3315 (n2176, n1392, n_1780);
  not g3316 (n_1781, n2176);
  and g3317 (n2177, n1396, n_1781);
  not g3318 (n_1782, n2177);
  and g3319 (n2178, n1663, n_1782);
  not g3320 (n_1783, n2178);
  and g3321 (n2179, n392, n_1783);
  not g3322 (n_1784, n2179);
  and g3323 (n2180, n396, n_1784);
  not g3324 (n_1785, n2180);
  and g3325 (n2181, n400, n_1785);
  not g3326 (n_1786, n2181);
  and g3327 (n2182, n404, n_1786);
  not g3328 (n_1787, n2182);
  and g3329 (n2183, n408, n_1787);
  and g3330 (n2184, \req[11] , n_52);
  not g3331 (n_1788, n2183);
  and g3332 (\grant[11] , n_1788, n2184);
  not g3333 (n_1789, n754);
  and g3334 (n2186, n419, n_1789);
  not g3335 (n_1790, n2186);
  and g3336 (n2187, n424, n_1790);
  not g3337 (n_1791, n2187);
  and g3338 (n2188, n428, n_1791);
  not g3339 (n_1792, n2188);
  and g3340 (n2189, n432, n_1792);
  not g3341 (n_1793, n2189);
  and g3342 (n2190, n436, n_1793);
  not g3343 (n_1794, n2190);
  and g3344 (n2191, n440, n_1794);
  not g3345 (n_1795, n2191);
  and g3346 (n2192, n444, n_1795);
  not g3347 (n_1796, n2192);
  and g3348 (n2193, n448, n_1796);
  not g3349 (n_1797, n2193);
  and g3350 (n2194, n452, n_1797);
  not g3351 (n_1798, n2194);
  and g3352 (n2195, n456, n_1798);
  not g3353 (n_1799, n2195);
  and g3354 (n2196, n460, n_1799);
  not g3355 (n_1800, n2196);
  and g3356 (n2197, n464, n_1800);
  not g3357 (n_1801, n2197);
  and g3358 (n2198, n468, n_1801);
  not g3359 (n_1802, n2198);
  and g3360 (n2199, n472, n_1802);
  not g3361 (n_1803, n2199);
  and g3362 (n2200, n476, n_1803);
  not g3363 (n_1804, n2200);
  and g3364 (n2201, n480, n_1804);
  not g3365 (n_1805, n2201);
  and g3366 (n2202, n484, n_1805);
  not g3367 (n_1806, n2202);
  and g3368 (n2203, n488, n_1806);
  not g3369 (n_1807, n2203);
  and g3370 (n2204, n492, n_1807);
  not g3371 (n_1808, n2204);
  and g3372 (n2205, n496, n_1808);
  not g3373 (n_1809, n2205);
  and g3374 (n2206, n500, n_1809);
  not g3375 (n_1810, n2206);
  and g3376 (n2207, n504, n_1810);
  not g3377 (n_1811, n2207);
  and g3378 (n2208, n508, n_1811);
  not g3379 (n_1812, n2208);
  and g3380 (n2209, n512, n_1812);
  not g3381 (n_1813, n2209);
  and g3382 (n2210, n516, n_1813);
  not g3383 (n_1814, n2210);
  and g3384 (n2211, n520, n_1814);
  not g3385 (n_1815, n2211);
  and g3386 (n2212, n524, n_1815);
  not g3387 (n_1816, n2212);
  and g3388 (n2213, n528, n_1816);
  not g3389 (n_1817, n2213);
  and g3390 (n2214, n532, n_1817);
  not g3391 (n_1818, n2214);
  and g3392 (n2215, n536, n_1818);
  not g3393 (n_1819, n2215);
  and g3394 (n2216, n540, n_1819);
  not g3395 (n_1820, n2216);
  and g3396 (n2217, n544, n_1820);
  not g3397 (n_1821, n2217);
  and g3398 (n2218, n548, n_1821);
  not g3399 (n_1822, n2218);
  and g3400 (n2219, n552, n_1822);
  not g3401 (n_1823, n2219);
  and g3402 (n2220, n556, n_1823);
  not g3403 (n_1824, n2220);
  and g3404 (n2221, n560, n_1824);
  not g3405 (n_1825, n2221);
  and g3406 (n2222, n564, n_1825);
  not g3407 (n_1826, n2222);
  and g3408 (n2223, n568, n_1826);
  not g3409 (n_1827, n2223);
  and g3410 (n2224, n572, n_1827);
  not g3411 (n_1828, n2224);
  and g3412 (n2225, n576, n_1828);
  not g3413 (n_1829, n2225);
  and g3414 (n2226, n580, n_1829);
  not g3415 (n_1830, n2226);
  and g3416 (n2227, n584, n_1830);
  not g3417 (n_1831, n2227);
  and g3418 (n2228, n588, n_1831);
  not g3419 (n_1832, n2228);
  and g3420 (n2229, n592, n_1832);
  not g3421 (n_1833, n2229);
  and g3422 (n2230, n596, n_1833);
  not g3423 (n_1834, n2230);
  and g3424 (n2231, n600, n_1834);
  not g3425 (n_1835, n2231);
  and g3426 (n2232, n604, n_1835);
  not g3427 (n_1836, n2232);
  and g3428 (n2233, n608, n_1836);
  not g3429 (n_1837, n2233);
  and g3430 (n2234, n612, n_1837);
  not g3431 (n_1838, n2234);
  and g3432 (n2235, n616, n_1838);
  not g3433 (n_1839, n2235);
  and g3434 (n2236, n620, n_1839);
  not g3435 (n_1840, n2236);
  and g3436 (n2237, n624, n_1840);
  not g3437 (n_1841, n2237);
  and g3438 (n2238, n628, n_1841);
  not g3439 (n_1842, n2238);
  and g3440 (n2239, n632, n_1842);
  not g3441 (n_1843, n2239);
  and g3442 (n2240, n636, n_1843);
  not g3443 (n_1844, n2240);
  and g3444 (n2241, n640, n_1844);
  not g3445 (n_1845, n2241);
  and g3446 (n2242, n644, n_1845);
  not g3447 (n_1846, n2242);
  and g3448 (n2243, n648, n_1846);
  not g3449 (n_1847, n2243);
  and g3450 (n2244, n652, n_1847);
  not g3451 (n_1848, n2244);
  and g3452 (n2245, n656, n_1848);
  not g3453 (n_1849, n2245);
  and g3454 (n2246, n660, n_1849);
  not g3455 (n_1850, n2246);
  and g3456 (n2247, n664, n_1850);
  not g3457 (n_1851, n2247);
  and g3458 (n2248, n668, n_1851);
  not g3459 (n_1852, n2248);
  and g3460 (n2249, n672, n_1852);
  not g3461 (n_1853, n2249);
  and g3462 (n2250, n676, n_1853);
  not g3463 (n_1854, n2250);
  and g3464 (n2251, n680, n_1854);
  not g3465 (n_1855, n2251);
  and g3466 (n2252, n684, n_1855);
  not g3467 (n_1856, n2252);
  and g3468 (n2253, n688, n_1856);
  not g3469 (n_1857, n2253);
  and g3470 (n2254, n692, n_1857);
  not g3471 (n_1858, n2254);
  and g3472 (n2255, n696, n_1858);
  not g3473 (n_1859, n2255);
  and g3474 (n2256, n700, n_1859);
  not g3475 (n_1860, n2256);
  and g3476 (n2257, n704, n_1860);
  not g3477 (n_1861, n2257);
  and g3478 (n2258, n708, n_1861);
  not g3479 (n_1862, n2258);
  and g3480 (n2259, n712, n_1862);
  not g3481 (n_1863, n2259);
  and g3482 (n2260, n716, n_1863);
  not g3483 (n_1864, n2260);
  and g3484 (n2261, n720, n_1864);
  not g3485 (n_1865, n2261);
  and g3486 (n2262, n1484, n_1865);
  not g3487 (n_1866, n2262);
  and g3488 (n2263, n1486, n_1866);
  not g3489 (n_1867, n2263);
  and g3490 (n2264, n1750, n_1867);
  not g3491 (n_1868, n2264);
  and g3492 (n2265, n731, n_1868);
  not g3493 (n_1869, n2265);
  and g3494 (n2266, n735, n_1869);
  not g3495 (n_1870, n2266);
  and g3496 (n2267, n739, n_1870);
  not g3497 (n_1871, n2267);
  and g3498 (n2268, n743, n_1871);
  not g3499 (n_1872, n2268);
  and g3500 (n2269, n747, n_1872);
  and g3501 (n2270, \req[12] , n_617);
  not g3502 (n_1873, n2269);
  and g3503 (\grant[12] , n_1873, n2270);
  not g3504 (n_1874, n1091);
  and g3505 (n2272, n758, n_1874);
  not g3506 (n_1875, n2272);
  and g3507 (n2273, n763, n_1875);
  not g3508 (n_1876, n2273);
  and g3509 (n2274, n767, n_1876);
  not g3510 (n_1877, n2274);
  and g3511 (n2275, n771, n_1877);
  not g3512 (n_1878, n2275);
  and g3513 (n2276, n775, n_1878);
  not g3514 (n_1879, n2276);
  and g3515 (n2277, n779, n_1879);
  not g3516 (n_1880, n2277);
  and g3517 (n2278, n783, n_1880);
  not g3518 (n_1881, n2278);
  and g3519 (n2279, n787, n_1881);
  not g3520 (n_1882, n2279);
  and g3521 (n2280, n791, n_1882);
  not g3522 (n_1883, n2280);
  and g3523 (n2281, n795, n_1883);
  not g3524 (n_1884, n2281);
  and g3525 (n2282, n799, n_1884);
  not g3526 (n_1885, n2282);
  and g3527 (n2283, n803, n_1885);
  not g3528 (n_1886, n2283);
  and g3529 (n2284, n807, n_1886);
  not g3530 (n_1887, n2284);
  and g3531 (n2285, n811, n_1887);
  not g3532 (n_1888, n2285);
  and g3533 (n2286, n815, n_1888);
  not g3534 (n_1889, n2286);
  and g3535 (n2287, n819, n_1889);
  not g3536 (n_1890, n2287);
  and g3537 (n2288, n823, n_1890);
  not g3538 (n_1891, n2288);
  and g3539 (n2289, n827, n_1891);
  not g3540 (n_1892, n2289);
  and g3541 (n2290, n831, n_1892);
  not g3542 (n_1893, n2290);
  and g3543 (n2291, n835, n_1893);
  not g3544 (n_1894, n2291);
  and g3545 (n2292, n839, n_1894);
  not g3546 (n_1895, n2292);
  and g3547 (n2293, n843, n_1895);
  not g3548 (n_1896, n2293);
  and g3549 (n2294, n847, n_1896);
  not g3550 (n_1897, n2294);
  and g3551 (n2295, n851, n_1897);
  not g3552 (n_1898, n2295);
  and g3553 (n2296, n855, n_1898);
  not g3554 (n_1899, n2296);
  and g3555 (n2297, n859, n_1899);
  not g3556 (n_1900, n2297);
  and g3557 (n2298, n863, n_1900);
  not g3558 (n_1901, n2298);
  and g3559 (n2299, n867, n_1901);
  not g3560 (n_1902, n2299);
  and g3561 (n2300, n871, n_1902);
  not g3562 (n_1903, n2300);
  and g3563 (n2301, n875, n_1903);
  not g3564 (n_1904, n2301);
  and g3565 (n2302, n879, n_1904);
  not g3566 (n_1905, n2302);
  and g3567 (n2303, n883, n_1905);
  not g3568 (n_1906, n2303);
  and g3569 (n2304, n887, n_1906);
  not g3570 (n_1907, n2304);
  and g3571 (n2305, n891, n_1907);
  not g3572 (n_1908, n2305);
  and g3573 (n2306, n895, n_1908);
  not g3574 (n_1909, n2306);
  and g3575 (n2307, n899, n_1909);
  not g3576 (n_1910, n2307);
  and g3577 (n2308, n903, n_1910);
  not g3578 (n_1911, n2308);
  and g3579 (n2309, n907, n_1911);
  not g3580 (n_1912, n2309);
  and g3581 (n2310, n911, n_1912);
  not g3582 (n_1913, n2310);
  and g3583 (n2311, n915, n_1913);
  not g3584 (n_1914, n2311);
  and g3585 (n2312, n919, n_1914);
  not g3586 (n_1915, n2312);
  and g3587 (n2313, n923, n_1915);
  not g3588 (n_1916, n2313);
  and g3589 (n2314, n927, n_1916);
  not g3590 (n_1917, n2314);
  and g3591 (n2315, n931, n_1917);
  not g3592 (n_1918, n2315);
  and g3593 (n2316, n935, n_1918);
  not g3594 (n_1919, n2316);
  and g3595 (n2317, n939, n_1919);
  not g3596 (n_1920, n2317);
  and g3597 (n2318, n943, n_1920);
  not g3598 (n_1921, n2318);
  and g3599 (n2319, n947, n_1921);
  not g3600 (n_1922, n2319);
  and g3601 (n2320, n951, n_1922);
  not g3602 (n_1923, n2320);
  and g3603 (n2321, n955, n_1923);
  not g3604 (n_1924, n2321);
  and g3605 (n2322, n959, n_1924);
  not g3606 (n_1925, n2322);
  and g3607 (n2323, n963, n_1925);
  not g3608 (n_1926, n2323);
  and g3609 (n2324, n967, n_1926);
  not g3610 (n_1927, n2324);
  and g3611 (n2325, n971, n_1927);
  not g3612 (n_1928, n2325);
  and g3613 (n2326, n975, n_1928);
  not g3614 (n_1929, n2326);
  and g3615 (n2327, n979, n_1929);
  not g3616 (n_1930, n2327);
  and g3617 (n2328, n983, n_1930);
  not g3618 (n_1931, n2328);
  and g3619 (n2329, n987, n_1931);
  not g3620 (n_1932, n2329);
  and g3621 (n2330, n991, n_1932);
  not g3622 (n_1933, n2330);
  and g3623 (n2331, n995, n_1933);
  not g3624 (n_1934, n2331);
  and g3625 (n2332, n999, n_1934);
  not g3626 (n_1935, n2332);
  and g3627 (n2333, n1003, n_1935);
  not g3628 (n_1936, n2333);
  and g3629 (n2334, n1007, n_1936);
  not g3630 (n_1937, n2334);
  and g3631 (n2335, n1011, n_1937);
  not g3632 (n_1938, n2335);
  and g3633 (n2336, n1015, n_1938);
  not g3634 (n_1939, n2336);
  and g3635 (n2337, n1019, n_1939);
  not g3636 (n_1940, n2337);
  and g3637 (n2338, n1023, n_1940);
  not g3638 (n_1941, n2338);
  and g3639 (n2339, n1027, n_1941);
  not g3640 (n_1942, n2339);
  and g3641 (n2340, n1031, n_1942);
  not g3642 (n_1943, n2340);
  and g3643 (n2341, n1035, n_1943);
  not g3644 (n_1944, n2341);
  and g3645 (n2342, n1039, n_1944);
  not g3646 (n_1945, n2342);
  and g3647 (n2343, n1043, n_1945);
  not g3648 (n_1946, n2343);
  and g3649 (n2344, n1047, n_1946);
  not g3650 (n_1947, n2344);
  and g3651 (n2345, n1051, n_1947);
  not g3652 (n_1948, n2345);
  and g3653 (n2346, n1055, n_1948);
  not g3654 (n_1949, n2346);
  and g3655 (n2347, n1059, n_1949);
  not g3656 (n_1950, n2347);
  and g3657 (n2348, n1574, n_1950);
  not g3658 (n_1951, n2348);
  and g3659 (n2349, n1576, n_1951);
  not g3660 (n_1952, n2349);
  and g3661 (n2350, n1837, n_1952);
  not g3662 (n_1953, n2350);
  and g3663 (n2351, n1068, n_1953);
  not g3664 (n_1954, n2351);
  and g3665 (n2352, n1072, n_1954);
  not g3666 (n_1955, n2352);
  and g3667 (n2353, n1076, n_1955);
  not g3668 (n_1956, n2353);
  and g3669 (n2354, n1080, n_1956);
  not g3670 (n_1957, n2354);
  and g3671 (n2355, n1084, n_1957);
  and g3672 (n2356, \req[13] , n_863);
  not g3673 (n_1958, n2355);
  and g3674 (\grant[13] , n_1958, n2356);
  not g3675 (n_1959, n423);
  and g3676 (n2358, n_1959, n1095);
  not g3677 (n_1960, n2358);
  and g3678 (n2359, n1100, n_1960);
  not g3679 (n_1961, n2359);
  and g3680 (n2360, n1104, n_1961);
  not g3681 (n_1962, n2360);
  and g3682 (n2361, n1108, n_1962);
  not g3683 (n_1963, n2361);
  and g3684 (n2362, n1112, n_1963);
  not g3685 (n_1964, n2362);
  and g3686 (n2363, n1116, n_1964);
  not g3687 (n_1965, n2363);
  and g3688 (n2364, n1120, n_1965);
  not g3689 (n_1966, n2364);
  and g3690 (n2365, n1124, n_1966);
  not g3691 (n_1967, n2365);
  and g3692 (n2366, n1128, n_1967);
  not g3693 (n_1968, n2366);
  and g3694 (n2367, n1132, n_1968);
  not g3695 (n_1969, n2367);
  and g3696 (n2368, n1136, n_1969);
  not g3697 (n_1970, n2368);
  and g3698 (n2369, n1140, n_1970);
  not g3699 (n_1971, n2369);
  and g3700 (n2370, n1144, n_1971);
  not g3701 (n_1972, n2370);
  and g3702 (n2371, n1148, n_1972);
  not g3703 (n_1973, n2371);
  and g3704 (n2372, n1152, n_1973);
  not g3705 (n_1974, n2372);
  and g3706 (n2373, n1156, n_1974);
  not g3707 (n_1975, n2373);
  and g3708 (n2374, n1160, n_1975);
  not g3709 (n_1976, n2374);
  and g3710 (n2375, n1164, n_1976);
  not g3711 (n_1977, n2375);
  and g3712 (n2376, n1168, n_1977);
  not g3713 (n_1978, n2376);
  and g3714 (n2377, n1172, n_1978);
  not g3715 (n_1979, n2377);
  and g3716 (n2378, n1176, n_1979);
  not g3717 (n_1980, n2378);
  and g3718 (n2379, n1180, n_1980);
  not g3719 (n_1981, n2379);
  and g3720 (n2380, n1184, n_1981);
  not g3721 (n_1982, n2380);
  and g3722 (n2381, n1188, n_1982);
  not g3723 (n_1983, n2381);
  and g3724 (n2382, n1192, n_1983);
  not g3725 (n_1984, n2382);
  and g3726 (n2383, n1196, n_1984);
  not g3727 (n_1985, n2383);
  and g3728 (n2384, n1200, n_1985);
  not g3729 (n_1986, n2384);
  and g3730 (n2385, n1204, n_1986);
  not g3731 (n_1987, n2385);
  and g3732 (n2386, n1208, n_1987);
  not g3733 (n_1988, n2386);
  and g3734 (n2387, n1212, n_1988);
  not g3735 (n_1989, n2387);
  and g3736 (n2388, n1216, n_1989);
  not g3737 (n_1990, n2388);
  and g3738 (n2389, n1220, n_1990);
  not g3739 (n_1991, n2389);
  and g3740 (n2390, n1224, n_1991);
  not g3741 (n_1992, n2390);
  and g3742 (n2391, n1228, n_1992);
  not g3743 (n_1993, n2391);
  and g3744 (n2392, n1232, n_1993);
  not g3745 (n_1994, n2392);
  and g3746 (n2393, n1236, n_1994);
  not g3747 (n_1995, n2393);
  and g3748 (n2394, n1240, n_1995);
  not g3749 (n_1996, n2394);
  and g3750 (n2395, n1244, n_1996);
  not g3751 (n_1997, n2395);
  and g3752 (n2396, n1248, n_1997);
  not g3753 (n_1998, n2396);
  and g3754 (n2397, n1252, n_1998);
  not g3755 (n_1999, n2397);
  and g3756 (n2398, n1256, n_1999);
  not g3757 (n_2000, n2398);
  and g3758 (n2399, n1260, n_2000);
  not g3759 (n_2001, n2399);
  and g3760 (n2400, n1264, n_2001);
  not g3761 (n_2002, n2400);
  and g3762 (n2401, n1268, n_2002);
  not g3763 (n_2003, n2401);
  and g3764 (n2402, n1272, n_2003);
  not g3765 (n_2004, n2402);
  and g3766 (n2403, n1276, n_2004);
  not g3767 (n_2005, n2403);
  and g3768 (n2404, n1280, n_2005);
  not g3769 (n_2006, n2404);
  and g3770 (n2405, n1284, n_2006);
  not g3771 (n_2007, n2405);
  and g3772 (n2406, n1288, n_2007);
  not g3773 (n_2008, n2406);
  and g3774 (n2407, n1292, n_2008);
  not g3775 (n_2009, n2407);
  and g3776 (n2408, n1296, n_2009);
  not g3777 (n_2010, n2408);
  and g3778 (n2409, n1300, n_2010);
  not g3779 (n_2011, n2409);
  and g3780 (n2410, n1304, n_2011);
  not g3781 (n_2012, n2410);
  and g3782 (n2411, n1308, n_2012);
  not g3783 (n_2013, n2411);
  and g3784 (n2412, n1312, n_2013);
  not g3785 (n_2014, n2412);
  and g3786 (n2413, n1316, n_2014);
  not g3787 (n_2015, n2413);
  and g3788 (n2414, n1320, n_2015);
  not g3789 (n_2016, n2414);
  and g3790 (n2415, n1324, n_2016);
  not g3791 (n_2017, n2415);
  and g3792 (n2416, n1328, n_2017);
  not g3793 (n_2018, n2416);
  and g3794 (n2417, n1332, n_2018);
  not g3795 (n_2019, n2417);
  and g3796 (n2418, n1336, n_2019);
  not g3797 (n_2020, n2418);
  and g3798 (n2419, n1340, n_2020);
  not g3799 (n_2021, n2419);
  and g3800 (n2420, n1344, n_2021);
  not g3801 (n_2022, n2420);
  and g3802 (n2421, n1348, n_2022);
  not g3803 (n_2023, n2421);
  and g3804 (n2422, n1352, n_2023);
  not g3805 (n_2024, n2422);
  and g3806 (n2423, n1356, n_2024);
  not g3807 (n_2025, n2423);
  and g3808 (n2424, n1360, n_2025);
  not g3809 (n_2026, n2424);
  and g3810 (n2425, n1364, n_2026);
  not g3811 (n_2027, n2425);
  and g3812 (n2426, n1368, n_2027);
  not g3813 (n_2028, n2426);
  and g3814 (n2427, n1372, n_2028);
  not g3815 (n_2029, n2427);
  and g3816 (n2428, n1376, n_2029);
  not g3817 (n_2030, n2428);
  and g3818 (n2429, n1380, n_2030);
  not g3819 (n_2031, n2429);
  and g3820 (n2430, n1384, n_2031);
  not g3821 (n_2032, n2430);
  and g3822 (n2431, n1388, n_2032);
  not g3823 (n_2033, n2431);
  and g3824 (n2432, n1392, n_2033);
  not g3825 (n_2034, n2432);
  and g3826 (n2433, n1396, n_2034);
  not g3827 (n_2035, n2433);
  and g3828 (n2434, n1663, n_2035);
  not g3829 (n_2036, n2434);
  and g3830 (n2435, n392, n_2036);
  not g3831 (n_2037, n2435);
  and g3832 (n2436, n396, n_2037);
  not g3833 (n_2038, n2436);
  and g3834 (n2437, n400, n_2038);
  not g3835 (n_2039, n2437);
  and g3836 (n2438, n404, n_2039);
  not g3837 (n_2040, n2438);
  and g3838 (n2439, n408, n_2040);
  not g3839 (n_2041, n2439);
  and g3840 (n2440, n412, n_2041);
  not g3841 (n_2042, n2440);
  and g3842 (n2441, n416, n_2042);
  and g3843 (n2442, \req[14] , n_66);
  not g3844 (n_2043, n2441);
  and g3845 (\grant[14] , n_2043, n2442);
  not g3846 (n_2044, n762);
  and g3847 (n2444, n427, n_2044);
  not g3848 (n_2045, n2444);
  and g3849 (n2445, n432, n_2045);
  not g3850 (n_2046, n2445);
  and g3851 (n2446, n436, n_2046);
  not g3852 (n_2047, n2446);
  and g3853 (n2447, n440, n_2047);
  not g3854 (n_2048, n2447);
  and g3855 (n2448, n444, n_2048);
  not g3856 (n_2049, n2448);
  and g3857 (n2449, n448, n_2049);
  not g3858 (n_2050, n2449);
  and g3859 (n2450, n452, n_2050);
  not g3860 (n_2051, n2450);
  and g3861 (n2451, n456, n_2051);
  not g3862 (n_2052, n2451);
  and g3863 (n2452, n460, n_2052);
  not g3864 (n_2053, n2452);
  and g3865 (n2453, n464, n_2053);
  not g3866 (n_2054, n2453);
  and g3867 (n2454, n468, n_2054);
  not g3868 (n_2055, n2454);
  and g3869 (n2455, n472, n_2055);
  not g3870 (n_2056, n2455);
  and g3871 (n2456, n476, n_2056);
  not g3872 (n_2057, n2456);
  and g3873 (n2457, n480, n_2057);
  not g3874 (n_2058, n2457);
  and g3875 (n2458, n484, n_2058);
  not g3876 (n_2059, n2458);
  and g3877 (n2459, n488, n_2059);
  not g3878 (n_2060, n2459);
  and g3879 (n2460, n492, n_2060);
  not g3880 (n_2061, n2460);
  and g3881 (n2461, n496, n_2061);
  not g3882 (n_2062, n2461);
  and g3883 (n2462, n500, n_2062);
  not g3884 (n_2063, n2462);
  and g3885 (n2463, n504, n_2063);
  not g3886 (n_2064, n2463);
  and g3887 (n2464, n508, n_2064);
  not g3888 (n_2065, n2464);
  and g3889 (n2465, n512, n_2065);
  not g3890 (n_2066, n2465);
  and g3891 (n2466, n516, n_2066);
  not g3892 (n_2067, n2466);
  and g3893 (n2467, n520, n_2067);
  not g3894 (n_2068, n2467);
  and g3895 (n2468, n524, n_2068);
  not g3896 (n_2069, n2468);
  and g3897 (n2469, n528, n_2069);
  not g3898 (n_2070, n2469);
  and g3899 (n2470, n532, n_2070);
  not g3900 (n_2071, n2470);
  and g3901 (n2471, n536, n_2071);
  not g3902 (n_2072, n2471);
  and g3903 (n2472, n540, n_2072);
  not g3904 (n_2073, n2472);
  and g3905 (n2473, n544, n_2073);
  not g3906 (n_2074, n2473);
  and g3907 (n2474, n548, n_2074);
  not g3908 (n_2075, n2474);
  and g3909 (n2475, n552, n_2075);
  not g3910 (n_2076, n2475);
  and g3911 (n2476, n556, n_2076);
  not g3912 (n_2077, n2476);
  and g3913 (n2477, n560, n_2077);
  not g3914 (n_2078, n2477);
  and g3915 (n2478, n564, n_2078);
  not g3916 (n_2079, n2478);
  and g3917 (n2479, n568, n_2079);
  not g3918 (n_2080, n2479);
  and g3919 (n2480, n572, n_2080);
  not g3920 (n_2081, n2480);
  and g3921 (n2481, n576, n_2081);
  not g3922 (n_2082, n2481);
  and g3923 (n2482, n580, n_2082);
  not g3924 (n_2083, n2482);
  and g3925 (n2483, n584, n_2083);
  not g3926 (n_2084, n2483);
  and g3927 (n2484, n588, n_2084);
  not g3928 (n_2085, n2484);
  and g3929 (n2485, n592, n_2085);
  not g3930 (n_2086, n2485);
  and g3931 (n2486, n596, n_2086);
  not g3932 (n_2087, n2486);
  and g3933 (n2487, n600, n_2087);
  not g3934 (n_2088, n2487);
  and g3935 (n2488, n604, n_2088);
  not g3936 (n_2089, n2488);
  and g3937 (n2489, n608, n_2089);
  not g3938 (n_2090, n2489);
  and g3939 (n2490, n612, n_2090);
  not g3940 (n_2091, n2490);
  and g3941 (n2491, n616, n_2091);
  not g3942 (n_2092, n2491);
  and g3943 (n2492, n620, n_2092);
  not g3944 (n_2093, n2492);
  and g3945 (n2493, n624, n_2093);
  not g3946 (n_2094, n2493);
  and g3947 (n2494, n628, n_2094);
  not g3948 (n_2095, n2494);
  and g3949 (n2495, n632, n_2095);
  not g3950 (n_2096, n2495);
  and g3951 (n2496, n636, n_2096);
  not g3952 (n_2097, n2496);
  and g3953 (n2497, n640, n_2097);
  not g3954 (n_2098, n2497);
  and g3955 (n2498, n644, n_2098);
  not g3956 (n_2099, n2498);
  and g3957 (n2499, n648, n_2099);
  not g3958 (n_2100, n2499);
  and g3959 (n2500, n652, n_2100);
  not g3960 (n_2101, n2500);
  and g3961 (n2501, n656, n_2101);
  not g3962 (n_2102, n2501);
  and g3963 (n2502, n660, n_2102);
  not g3964 (n_2103, n2502);
  and g3965 (n2503, n664, n_2103);
  not g3966 (n_2104, n2503);
  and g3967 (n2504, n668, n_2104);
  not g3968 (n_2105, n2504);
  and g3969 (n2505, n672, n_2105);
  not g3970 (n_2106, n2505);
  and g3971 (n2506, n676, n_2106);
  not g3972 (n_2107, n2506);
  and g3973 (n2507, n680, n_2107);
  not g3974 (n_2108, n2507);
  and g3975 (n2508, n684, n_2108);
  not g3976 (n_2109, n2508);
  and g3977 (n2509, n688, n_2109);
  not g3978 (n_2110, n2509);
  and g3979 (n2510, n692, n_2110);
  not g3980 (n_2111, n2510);
  and g3981 (n2511, n696, n_2111);
  not g3982 (n_2112, n2511);
  and g3983 (n2512, n700, n_2112);
  not g3984 (n_2113, n2512);
  and g3985 (n2513, n704, n_2113);
  not g3986 (n_2114, n2513);
  and g3987 (n2514, n708, n_2114);
  not g3988 (n_2115, n2514);
  and g3989 (n2515, n712, n_2115);
  not g3990 (n_2116, n2515);
  and g3991 (n2516, n716, n_2116);
  not g3992 (n_2117, n2516);
  and g3993 (n2517, n720, n_2117);
  not g3994 (n_2118, n2517);
  and g3995 (n2518, n1484, n_2118);
  not g3996 (n_2119, n2518);
  and g3997 (n2519, n1486, n_2119);
  not g3998 (n_2120, n2519);
  and g3999 (n2520, n1750, n_2120);
  not g4000 (n_2121, n2520);
  and g4001 (n2521, n731, n_2121);
  not g4002 (n_2122, n2521);
  and g4003 (n2522, n735, n_2122);
  not g4004 (n_2123, n2522);
  and g4005 (n2523, n739, n_2123);
  not g4006 (n_2124, n2523);
  and g4007 (n2524, n743, n_2124);
  not g4008 (n_2125, n2524);
  and g4009 (n2525, n747, n_2125);
  not g4010 (n_2126, n2525);
  and g4011 (n2526, n751, n_2126);
  not g4012 (n_2127, n2526);
  and g4013 (n2527, n755, n_2127);
  and g4014 (n2528, \req[15] , n_623);
  not g4015 (n_2128, n2527);
  and g4016 (\grant[15] , n_2128, n2528);
  not g4017 (n_2129, n1099);
  and g4018 (n2530, n766, n_2129);
  not g4019 (n_2130, n2530);
  and g4020 (n2531, n771, n_2130);
  not g4021 (n_2131, n2531);
  and g4022 (n2532, n775, n_2131);
  not g4023 (n_2132, n2532);
  and g4024 (n2533, n779, n_2132);
  not g4025 (n_2133, n2533);
  and g4026 (n2534, n783, n_2133);
  not g4027 (n_2134, n2534);
  and g4028 (n2535, n787, n_2134);
  not g4029 (n_2135, n2535);
  and g4030 (n2536, n791, n_2135);
  not g4031 (n_2136, n2536);
  and g4032 (n2537, n795, n_2136);
  not g4033 (n_2137, n2537);
  and g4034 (n2538, n799, n_2137);
  not g4035 (n_2138, n2538);
  and g4036 (n2539, n803, n_2138);
  not g4037 (n_2139, n2539);
  and g4038 (n2540, n807, n_2139);
  not g4039 (n_2140, n2540);
  and g4040 (n2541, n811, n_2140);
  not g4041 (n_2141, n2541);
  and g4042 (n2542, n815, n_2141);
  not g4043 (n_2142, n2542);
  and g4044 (n2543, n819, n_2142);
  not g4045 (n_2143, n2543);
  and g4046 (n2544, n823, n_2143);
  not g4047 (n_2144, n2544);
  and g4048 (n2545, n827, n_2144);
  not g4049 (n_2145, n2545);
  and g4050 (n2546, n831, n_2145);
  not g4051 (n_2146, n2546);
  and g4052 (n2547, n835, n_2146);
  not g4053 (n_2147, n2547);
  and g4054 (n2548, n839, n_2147);
  not g4055 (n_2148, n2548);
  and g4056 (n2549, n843, n_2148);
  not g4057 (n_2149, n2549);
  and g4058 (n2550, n847, n_2149);
  not g4059 (n_2150, n2550);
  and g4060 (n2551, n851, n_2150);
  not g4061 (n_2151, n2551);
  and g4062 (n2552, n855, n_2151);
  not g4063 (n_2152, n2552);
  and g4064 (n2553, n859, n_2152);
  not g4065 (n_2153, n2553);
  and g4066 (n2554, n863, n_2153);
  not g4067 (n_2154, n2554);
  and g4068 (n2555, n867, n_2154);
  not g4069 (n_2155, n2555);
  and g4070 (n2556, n871, n_2155);
  not g4071 (n_2156, n2556);
  and g4072 (n2557, n875, n_2156);
  not g4073 (n_2157, n2557);
  and g4074 (n2558, n879, n_2157);
  not g4075 (n_2158, n2558);
  and g4076 (n2559, n883, n_2158);
  not g4077 (n_2159, n2559);
  and g4078 (n2560, n887, n_2159);
  not g4079 (n_2160, n2560);
  and g4080 (n2561, n891, n_2160);
  not g4081 (n_2161, n2561);
  and g4082 (n2562, n895, n_2161);
  not g4083 (n_2162, n2562);
  and g4084 (n2563, n899, n_2162);
  not g4085 (n_2163, n2563);
  and g4086 (n2564, n903, n_2163);
  not g4087 (n_2164, n2564);
  and g4088 (n2565, n907, n_2164);
  not g4089 (n_2165, n2565);
  and g4090 (n2566, n911, n_2165);
  not g4091 (n_2166, n2566);
  and g4092 (n2567, n915, n_2166);
  not g4093 (n_2167, n2567);
  and g4094 (n2568, n919, n_2167);
  not g4095 (n_2168, n2568);
  and g4096 (n2569, n923, n_2168);
  not g4097 (n_2169, n2569);
  and g4098 (n2570, n927, n_2169);
  not g4099 (n_2170, n2570);
  and g4100 (n2571, n931, n_2170);
  not g4101 (n_2171, n2571);
  and g4102 (n2572, n935, n_2171);
  not g4103 (n_2172, n2572);
  and g4104 (n2573, n939, n_2172);
  not g4105 (n_2173, n2573);
  and g4106 (n2574, n943, n_2173);
  not g4107 (n_2174, n2574);
  and g4108 (n2575, n947, n_2174);
  not g4109 (n_2175, n2575);
  and g4110 (n2576, n951, n_2175);
  not g4111 (n_2176, n2576);
  and g4112 (n2577, n955, n_2176);
  not g4113 (n_2177, n2577);
  and g4114 (n2578, n959, n_2177);
  not g4115 (n_2178, n2578);
  and g4116 (n2579, n963, n_2178);
  not g4117 (n_2179, n2579);
  and g4118 (n2580, n967, n_2179);
  not g4119 (n_2180, n2580);
  and g4120 (n2581, n971, n_2180);
  not g4121 (n_2181, n2581);
  and g4122 (n2582, n975, n_2181);
  not g4123 (n_2182, n2582);
  and g4124 (n2583, n979, n_2182);
  not g4125 (n_2183, n2583);
  and g4126 (n2584, n983, n_2183);
  not g4127 (n_2184, n2584);
  and g4128 (n2585, n987, n_2184);
  not g4129 (n_2185, n2585);
  and g4130 (n2586, n991, n_2185);
  not g4131 (n_2186, n2586);
  and g4132 (n2587, n995, n_2186);
  not g4133 (n_2187, n2587);
  and g4134 (n2588, n999, n_2187);
  not g4135 (n_2188, n2588);
  and g4136 (n2589, n1003, n_2188);
  not g4137 (n_2189, n2589);
  and g4138 (n2590, n1007, n_2189);
  not g4139 (n_2190, n2590);
  and g4140 (n2591, n1011, n_2190);
  not g4141 (n_2191, n2591);
  and g4142 (n2592, n1015, n_2191);
  not g4143 (n_2192, n2592);
  and g4144 (n2593, n1019, n_2192);
  not g4145 (n_2193, n2593);
  and g4146 (n2594, n1023, n_2193);
  not g4147 (n_2194, n2594);
  and g4148 (n2595, n1027, n_2194);
  not g4149 (n_2195, n2595);
  and g4150 (n2596, n1031, n_2195);
  not g4151 (n_2196, n2596);
  and g4152 (n2597, n1035, n_2196);
  not g4153 (n_2197, n2597);
  and g4154 (n2598, n1039, n_2197);
  not g4155 (n_2198, n2598);
  and g4156 (n2599, n1043, n_2198);
  not g4157 (n_2199, n2599);
  and g4158 (n2600, n1047, n_2199);
  not g4159 (n_2200, n2600);
  and g4160 (n2601, n1051, n_2200);
  not g4161 (n_2201, n2601);
  and g4162 (n2602, n1055, n_2201);
  not g4163 (n_2202, n2602);
  and g4164 (n2603, n1059, n_2202);
  not g4165 (n_2203, n2603);
  and g4166 (n2604, n1574, n_2203);
  not g4167 (n_2204, n2604);
  and g4168 (n2605, n1576, n_2204);
  not g4169 (n_2205, n2605);
  and g4170 (n2606, n1837, n_2205);
  not g4171 (n_2206, n2606);
  and g4172 (n2607, n1068, n_2206);
  not g4173 (n_2207, n2607);
  and g4174 (n2608, n1072, n_2207);
  not g4175 (n_2208, n2608);
  and g4176 (n2609, n1076, n_2208);
  not g4177 (n_2209, n2609);
  and g4178 (n2610, n1080, n_2209);
  not g4179 (n_2210, n2610);
  and g4180 (n2611, n1084, n_2210);
  not g4181 (n_2211, n2611);
  and g4182 (n2612, n1088, n_2211);
  not g4183 (n_2212, n2612);
  and g4184 (n2613, n1092, n_2212);
  and g4185 (n2614, \req[16] , n_867);
  not g4186 (n_2213, n2613);
  and g4187 (\grant[16] , n_2213, n2614);
  not g4188 (n_2214, n431);
  and g4189 (n2616, n_2214, n1103);
  not g4190 (n_2215, n2616);
  and g4191 (n2617, n1108, n_2215);
  not g4192 (n_2216, n2617);
  and g4193 (n2618, n1112, n_2216);
  not g4194 (n_2217, n2618);
  and g4195 (n2619, n1116, n_2217);
  not g4196 (n_2218, n2619);
  and g4197 (n2620, n1120, n_2218);
  not g4198 (n_2219, n2620);
  and g4199 (n2621, n1124, n_2219);
  not g4200 (n_2220, n2621);
  and g4201 (n2622, n1128, n_2220);
  not g4202 (n_2221, n2622);
  and g4203 (n2623, n1132, n_2221);
  not g4204 (n_2222, n2623);
  and g4205 (n2624, n1136, n_2222);
  not g4206 (n_2223, n2624);
  and g4207 (n2625, n1140, n_2223);
  not g4208 (n_2224, n2625);
  and g4209 (n2626, n1144, n_2224);
  not g4210 (n_2225, n2626);
  and g4211 (n2627, n1148, n_2225);
  not g4212 (n_2226, n2627);
  and g4213 (n2628, n1152, n_2226);
  not g4214 (n_2227, n2628);
  and g4215 (n2629, n1156, n_2227);
  not g4216 (n_2228, n2629);
  and g4217 (n2630, n1160, n_2228);
  not g4218 (n_2229, n2630);
  and g4219 (n2631, n1164, n_2229);
  not g4220 (n_2230, n2631);
  and g4221 (n2632, n1168, n_2230);
  not g4222 (n_2231, n2632);
  and g4223 (n2633, n1172, n_2231);
  not g4224 (n_2232, n2633);
  and g4225 (n2634, n1176, n_2232);
  not g4226 (n_2233, n2634);
  and g4227 (n2635, n1180, n_2233);
  not g4228 (n_2234, n2635);
  and g4229 (n2636, n1184, n_2234);
  not g4230 (n_2235, n2636);
  and g4231 (n2637, n1188, n_2235);
  not g4232 (n_2236, n2637);
  and g4233 (n2638, n1192, n_2236);
  not g4234 (n_2237, n2638);
  and g4235 (n2639, n1196, n_2237);
  not g4236 (n_2238, n2639);
  and g4237 (n2640, n1200, n_2238);
  not g4238 (n_2239, n2640);
  and g4239 (n2641, n1204, n_2239);
  not g4240 (n_2240, n2641);
  and g4241 (n2642, n1208, n_2240);
  not g4242 (n_2241, n2642);
  and g4243 (n2643, n1212, n_2241);
  not g4244 (n_2242, n2643);
  and g4245 (n2644, n1216, n_2242);
  not g4246 (n_2243, n2644);
  and g4247 (n2645, n1220, n_2243);
  not g4248 (n_2244, n2645);
  and g4249 (n2646, n1224, n_2244);
  not g4250 (n_2245, n2646);
  and g4251 (n2647, n1228, n_2245);
  not g4252 (n_2246, n2647);
  and g4253 (n2648, n1232, n_2246);
  not g4254 (n_2247, n2648);
  and g4255 (n2649, n1236, n_2247);
  not g4256 (n_2248, n2649);
  and g4257 (n2650, n1240, n_2248);
  not g4258 (n_2249, n2650);
  and g4259 (n2651, n1244, n_2249);
  not g4260 (n_2250, n2651);
  and g4261 (n2652, n1248, n_2250);
  not g4262 (n_2251, n2652);
  and g4263 (n2653, n1252, n_2251);
  not g4264 (n_2252, n2653);
  and g4265 (n2654, n1256, n_2252);
  not g4266 (n_2253, n2654);
  and g4267 (n2655, n1260, n_2253);
  not g4268 (n_2254, n2655);
  and g4269 (n2656, n1264, n_2254);
  not g4270 (n_2255, n2656);
  and g4271 (n2657, n1268, n_2255);
  not g4272 (n_2256, n2657);
  and g4273 (n2658, n1272, n_2256);
  not g4274 (n_2257, n2658);
  and g4275 (n2659, n1276, n_2257);
  not g4276 (n_2258, n2659);
  and g4277 (n2660, n1280, n_2258);
  not g4278 (n_2259, n2660);
  and g4279 (n2661, n1284, n_2259);
  not g4280 (n_2260, n2661);
  and g4281 (n2662, n1288, n_2260);
  not g4282 (n_2261, n2662);
  and g4283 (n2663, n1292, n_2261);
  not g4284 (n_2262, n2663);
  and g4285 (n2664, n1296, n_2262);
  not g4286 (n_2263, n2664);
  and g4287 (n2665, n1300, n_2263);
  not g4288 (n_2264, n2665);
  and g4289 (n2666, n1304, n_2264);
  not g4290 (n_2265, n2666);
  and g4291 (n2667, n1308, n_2265);
  not g4292 (n_2266, n2667);
  and g4293 (n2668, n1312, n_2266);
  not g4294 (n_2267, n2668);
  and g4295 (n2669, n1316, n_2267);
  not g4296 (n_2268, n2669);
  and g4297 (n2670, n1320, n_2268);
  not g4298 (n_2269, n2670);
  and g4299 (n2671, n1324, n_2269);
  not g4300 (n_2270, n2671);
  and g4301 (n2672, n1328, n_2270);
  not g4302 (n_2271, n2672);
  and g4303 (n2673, n1332, n_2271);
  not g4304 (n_2272, n2673);
  and g4305 (n2674, n1336, n_2272);
  not g4306 (n_2273, n2674);
  and g4307 (n2675, n1340, n_2273);
  not g4308 (n_2274, n2675);
  and g4309 (n2676, n1344, n_2274);
  not g4310 (n_2275, n2676);
  and g4311 (n2677, n1348, n_2275);
  not g4312 (n_2276, n2677);
  and g4313 (n2678, n1352, n_2276);
  not g4314 (n_2277, n2678);
  and g4315 (n2679, n1356, n_2277);
  not g4316 (n_2278, n2679);
  and g4317 (n2680, n1360, n_2278);
  not g4318 (n_2279, n2680);
  and g4319 (n2681, n1364, n_2279);
  not g4320 (n_2280, n2681);
  and g4321 (n2682, n1368, n_2280);
  not g4322 (n_2281, n2682);
  and g4323 (n2683, n1372, n_2281);
  not g4324 (n_2282, n2683);
  and g4325 (n2684, n1376, n_2282);
  not g4326 (n_2283, n2684);
  and g4327 (n2685, n1380, n_2283);
  not g4328 (n_2284, n2685);
  and g4329 (n2686, n1384, n_2284);
  not g4330 (n_2285, n2686);
  and g4331 (n2687, n1388, n_2285);
  not g4332 (n_2286, n2687);
  and g4333 (n2688, n1392, n_2286);
  not g4334 (n_2287, n2688);
  and g4335 (n2689, n1396, n_2287);
  not g4336 (n_2288, n2689);
  and g4337 (n2690, n1663, n_2288);
  not g4338 (n_2289, n2690);
  and g4339 (n2691, n392, n_2289);
  not g4340 (n_2290, n2691);
  and g4341 (n2692, n396, n_2290);
  not g4342 (n_2291, n2692);
  and g4343 (n2693, n400, n_2291);
  not g4344 (n_2292, n2693);
  and g4345 (n2694, n404, n_2292);
  not g4346 (n_2293, n2694);
  and g4347 (n2695, n408, n_2293);
  not g4348 (n_2294, n2695);
  and g4349 (n2696, n412, n_2294);
  not g4350 (n_2295, n2696);
  and g4351 (n2697, n416, n_2295);
  not g4352 (n_2296, n2697);
  and g4353 (n2698, n420, n_2296);
  not g4354 (n_2297, n2698);
  and g4355 (n2699, n424, n_2297);
  and g4356 (n2700, \req[17] , n_80);
  not g4357 (n_2298, n2699);
  and g4358 (\grant[17] , n_2298, n2700);
  not g4359 (n_2299, n770);
  and g4360 (n2702, n435, n_2299);
  not g4361 (n_2300, n2702);
  and g4362 (n2703, n440, n_2300);
  not g4363 (n_2301, n2703);
  and g4364 (n2704, n444, n_2301);
  not g4365 (n_2302, n2704);
  and g4366 (n2705, n448, n_2302);
  not g4367 (n_2303, n2705);
  and g4368 (n2706, n452, n_2303);
  not g4369 (n_2304, n2706);
  and g4370 (n2707, n456, n_2304);
  not g4371 (n_2305, n2707);
  and g4372 (n2708, n460, n_2305);
  not g4373 (n_2306, n2708);
  and g4374 (n2709, n464, n_2306);
  not g4375 (n_2307, n2709);
  and g4376 (n2710, n468, n_2307);
  not g4377 (n_2308, n2710);
  and g4378 (n2711, n472, n_2308);
  not g4379 (n_2309, n2711);
  and g4380 (n2712, n476, n_2309);
  not g4381 (n_2310, n2712);
  and g4382 (n2713, n480, n_2310);
  not g4383 (n_2311, n2713);
  and g4384 (n2714, n484, n_2311);
  not g4385 (n_2312, n2714);
  and g4386 (n2715, n488, n_2312);
  not g4387 (n_2313, n2715);
  and g4388 (n2716, n492, n_2313);
  not g4389 (n_2314, n2716);
  and g4390 (n2717, n496, n_2314);
  not g4391 (n_2315, n2717);
  and g4392 (n2718, n500, n_2315);
  not g4393 (n_2316, n2718);
  and g4394 (n2719, n504, n_2316);
  not g4395 (n_2317, n2719);
  and g4396 (n2720, n508, n_2317);
  not g4397 (n_2318, n2720);
  and g4398 (n2721, n512, n_2318);
  not g4399 (n_2319, n2721);
  and g4400 (n2722, n516, n_2319);
  not g4401 (n_2320, n2722);
  and g4402 (n2723, n520, n_2320);
  not g4403 (n_2321, n2723);
  and g4404 (n2724, n524, n_2321);
  not g4405 (n_2322, n2724);
  and g4406 (n2725, n528, n_2322);
  not g4407 (n_2323, n2725);
  and g4408 (n2726, n532, n_2323);
  not g4409 (n_2324, n2726);
  and g4410 (n2727, n536, n_2324);
  not g4411 (n_2325, n2727);
  and g4412 (n2728, n540, n_2325);
  not g4413 (n_2326, n2728);
  and g4414 (n2729, n544, n_2326);
  not g4415 (n_2327, n2729);
  and g4416 (n2730, n548, n_2327);
  not g4417 (n_2328, n2730);
  and g4418 (n2731, n552, n_2328);
  not g4419 (n_2329, n2731);
  and g4420 (n2732, n556, n_2329);
  not g4421 (n_2330, n2732);
  and g4422 (n2733, n560, n_2330);
  not g4423 (n_2331, n2733);
  and g4424 (n2734, n564, n_2331);
  not g4425 (n_2332, n2734);
  and g4426 (n2735, n568, n_2332);
  not g4427 (n_2333, n2735);
  and g4428 (n2736, n572, n_2333);
  not g4429 (n_2334, n2736);
  and g4430 (n2737, n576, n_2334);
  not g4431 (n_2335, n2737);
  and g4432 (n2738, n580, n_2335);
  not g4433 (n_2336, n2738);
  and g4434 (n2739, n584, n_2336);
  not g4435 (n_2337, n2739);
  and g4436 (n2740, n588, n_2337);
  not g4437 (n_2338, n2740);
  and g4438 (n2741, n592, n_2338);
  not g4439 (n_2339, n2741);
  and g4440 (n2742, n596, n_2339);
  not g4441 (n_2340, n2742);
  and g4442 (n2743, n600, n_2340);
  not g4443 (n_2341, n2743);
  and g4444 (n2744, n604, n_2341);
  not g4445 (n_2342, n2744);
  and g4446 (n2745, n608, n_2342);
  not g4447 (n_2343, n2745);
  and g4448 (n2746, n612, n_2343);
  not g4449 (n_2344, n2746);
  and g4450 (n2747, n616, n_2344);
  not g4451 (n_2345, n2747);
  and g4452 (n2748, n620, n_2345);
  not g4453 (n_2346, n2748);
  and g4454 (n2749, n624, n_2346);
  not g4455 (n_2347, n2749);
  and g4456 (n2750, n628, n_2347);
  not g4457 (n_2348, n2750);
  and g4458 (n2751, n632, n_2348);
  not g4459 (n_2349, n2751);
  and g4460 (n2752, n636, n_2349);
  not g4461 (n_2350, n2752);
  and g4462 (n2753, n640, n_2350);
  not g4463 (n_2351, n2753);
  and g4464 (n2754, n644, n_2351);
  not g4465 (n_2352, n2754);
  and g4466 (n2755, n648, n_2352);
  not g4467 (n_2353, n2755);
  and g4468 (n2756, n652, n_2353);
  not g4469 (n_2354, n2756);
  and g4470 (n2757, n656, n_2354);
  not g4471 (n_2355, n2757);
  and g4472 (n2758, n660, n_2355);
  not g4473 (n_2356, n2758);
  and g4474 (n2759, n664, n_2356);
  not g4475 (n_2357, n2759);
  and g4476 (n2760, n668, n_2357);
  not g4477 (n_2358, n2760);
  and g4478 (n2761, n672, n_2358);
  not g4479 (n_2359, n2761);
  and g4480 (n2762, n676, n_2359);
  not g4481 (n_2360, n2762);
  and g4482 (n2763, n680, n_2360);
  not g4483 (n_2361, n2763);
  and g4484 (n2764, n684, n_2361);
  not g4485 (n_2362, n2764);
  and g4486 (n2765, n688, n_2362);
  not g4487 (n_2363, n2765);
  and g4488 (n2766, n692, n_2363);
  not g4489 (n_2364, n2766);
  and g4490 (n2767, n696, n_2364);
  not g4491 (n_2365, n2767);
  and g4492 (n2768, n700, n_2365);
  not g4493 (n_2366, n2768);
  and g4494 (n2769, n704, n_2366);
  not g4495 (n_2367, n2769);
  and g4496 (n2770, n708, n_2367);
  not g4497 (n_2368, n2770);
  and g4498 (n2771, n712, n_2368);
  not g4499 (n_2369, n2771);
  and g4500 (n2772, n716, n_2369);
  not g4501 (n_2370, n2772);
  and g4502 (n2773, n720, n_2370);
  not g4503 (n_2371, n2773);
  and g4504 (n2774, n1484, n_2371);
  not g4505 (n_2372, n2774);
  and g4506 (n2775, n1486, n_2372);
  not g4507 (n_2373, n2775);
  and g4508 (n2776, n1750, n_2373);
  not g4509 (n_2374, n2776);
  and g4510 (n2777, n731, n_2374);
  not g4511 (n_2375, n2777);
  and g4512 (n2778, n735, n_2375);
  not g4513 (n_2376, n2778);
  and g4514 (n2779, n739, n_2376);
  not g4515 (n_2377, n2779);
  and g4516 (n2780, n743, n_2377);
  not g4517 (n_2378, n2780);
  and g4518 (n2781, n747, n_2378);
  not g4519 (n_2379, n2781);
  and g4520 (n2782, n751, n_2379);
  not g4521 (n_2380, n2782);
  and g4522 (n2783, n755, n_2380);
  not g4523 (n_2381, n2783);
  and g4524 (n2784, n759, n_2381);
  not g4525 (n_2382, n2784);
  and g4526 (n2785, n763, n_2382);
  and g4527 (n2786, \req[18] , n_629);
  not g4528 (n_2383, n2785);
  and g4529 (\grant[18] , n_2383, n2786);
  not g4530 (n_2384, n1107);
  and g4531 (n2788, n774, n_2384);
  not g4532 (n_2385, n2788);
  and g4533 (n2789, n779, n_2385);
  not g4534 (n_2386, n2789);
  and g4535 (n2790, n783, n_2386);
  not g4536 (n_2387, n2790);
  and g4537 (n2791, n787, n_2387);
  not g4538 (n_2388, n2791);
  and g4539 (n2792, n791, n_2388);
  not g4540 (n_2389, n2792);
  and g4541 (n2793, n795, n_2389);
  not g4542 (n_2390, n2793);
  and g4543 (n2794, n799, n_2390);
  not g4544 (n_2391, n2794);
  and g4545 (n2795, n803, n_2391);
  not g4546 (n_2392, n2795);
  and g4547 (n2796, n807, n_2392);
  not g4548 (n_2393, n2796);
  and g4549 (n2797, n811, n_2393);
  not g4550 (n_2394, n2797);
  and g4551 (n2798, n815, n_2394);
  not g4552 (n_2395, n2798);
  and g4553 (n2799, n819, n_2395);
  not g4554 (n_2396, n2799);
  and g4555 (n2800, n823, n_2396);
  not g4556 (n_2397, n2800);
  and g4557 (n2801, n827, n_2397);
  not g4558 (n_2398, n2801);
  and g4559 (n2802, n831, n_2398);
  not g4560 (n_2399, n2802);
  and g4561 (n2803, n835, n_2399);
  not g4562 (n_2400, n2803);
  and g4563 (n2804, n839, n_2400);
  not g4564 (n_2401, n2804);
  and g4565 (n2805, n843, n_2401);
  not g4566 (n_2402, n2805);
  and g4567 (n2806, n847, n_2402);
  not g4568 (n_2403, n2806);
  and g4569 (n2807, n851, n_2403);
  not g4570 (n_2404, n2807);
  and g4571 (n2808, n855, n_2404);
  not g4572 (n_2405, n2808);
  and g4573 (n2809, n859, n_2405);
  not g4574 (n_2406, n2809);
  and g4575 (n2810, n863, n_2406);
  not g4576 (n_2407, n2810);
  and g4577 (n2811, n867, n_2407);
  not g4578 (n_2408, n2811);
  and g4579 (n2812, n871, n_2408);
  not g4580 (n_2409, n2812);
  and g4581 (n2813, n875, n_2409);
  not g4582 (n_2410, n2813);
  and g4583 (n2814, n879, n_2410);
  not g4584 (n_2411, n2814);
  and g4585 (n2815, n883, n_2411);
  not g4586 (n_2412, n2815);
  and g4587 (n2816, n887, n_2412);
  not g4588 (n_2413, n2816);
  and g4589 (n2817, n891, n_2413);
  not g4590 (n_2414, n2817);
  and g4591 (n2818, n895, n_2414);
  not g4592 (n_2415, n2818);
  and g4593 (n2819, n899, n_2415);
  not g4594 (n_2416, n2819);
  and g4595 (n2820, n903, n_2416);
  not g4596 (n_2417, n2820);
  and g4597 (n2821, n907, n_2417);
  not g4598 (n_2418, n2821);
  and g4599 (n2822, n911, n_2418);
  not g4600 (n_2419, n2822);
  and g4601 (n2823, n915, n_2419);
  not g4602 (n_2420, n2823);
  and g4603 (n2824, n919, n_2420);
  not g4604 (n_2421, n2824);
  and g4605 (n2825, n923, n_2421);
  not g4606 (n_2422, n2825);
  and g4607 (n2826, n927, n_2422);
  not g4608 (n_2423, n2826);
  and g4609 (n2827, n931, n_2423);
  not g4610 (n_2424, n2827);
  and g4611 (n2828, n935, n_2424);
  not g4612 (n_2425, n2828);
  and g4613 (n2829, n939, n_2425);
  not g4614 (n_2426, n2829);
  and g4615 (n2830, n943, n_2426);
  not g4616 (n_2427, n2830);
  and g4617 (n2831, n947, n_2427);
  not g4618 (n_2428, n2831);
  and g4619 (n2832, n951, n_2428);
  not g4620 (n_2429, n2832);
  and g4621 (n2833, n955, n_2429);
  not g4622 (n_2430, n2833);
  and g4623 (n2834, n959, n_2430);
  not g4624 (n_2431, n2834);
  and g4625 (n2835, n963, n_2431);
  not g4626 (n_2432, n2835);
  and g4627 (n2836, n967, n_2432);
  not g4628 (n_2433, n2836);
  and g4629 (n2837, n971, n_2433);
  not g4630 (n_2434, n2837);
  and g4631 (n2838, n975, n_2434);
  not g4632 (n_2435, n2838);
  and g4633 (n2839, n979, n_2435);
  not g4634 (n_2436, n2839);
  and g4635 (n2840, n983, n_2436);
  not g4636 (n_2437, n2840);
  and g4637 (n2841, n987, n_2437);
  not g4638 (n_2438, n2841);
  and g4639 (n2842, n991, n_2438);
  not g4640 (n_2439, n2842);
  and g4641 (n2843, n995, n_2439);
  not g4642 (n_2440, n2843);
  and g4643 (n2844, n999, n_2440);
  not g4644 (n_2441, n2844);
  and g4645 (n2845, n1003, n_2441);
  not g4646 (n_2442, n2845);
  and g4647 (n2846, n1007, n_2442);
  not g4648 (n_2443, n2846);
  and g4649 (n2847, n1011, n_2443);
  not g4650 (n_2444, n2847);
  and g4651 (n2848, n1015, n_2444);
  not g4652 (n_2445, n2848);
  and g4653 (n2849, n1019, n_2445);
  not g4654 (n_2446, n2849);
  and g4655 (n2850, n1023, n_2446);
  not g4656 (n_2447, n2850);
  and g4657 (n2851, n1027, n_2447);
  not g4658 (n_2448, n2851);
  and g4659 (n2852, n1031, n_2448);
  not g4660 (n_2449, n2852);
  and g4661 (n2853, n1035, n_2449);
  not g4662 (n_2450, n2853);
  and g4663 (n2854, n1039, n_2450);
  not g4664 (n_2451, n2854);
  and g4665 (n2855, n1043, n_2451);
  not g4666 (n_2452, n2855);
  and g4667 (n2856, n1047, n_2452);
  not g4668 (n_2453, n2856);
  and g4669 (n2857, n1051, n_2453);
  not g4670 (n_2454, n2857);
  and g4671 (n2858, n1055, n_2454);
  not g4672 (n_2455, n2858);
  and g4673 (n2859, n1059, n_2455);
  not g4674 (n_2456, n2859);
  and g4675 (n2860, n1574, n_2456);
  not g4676 (n_2457, n2860);
  and g4677 (n2861, n1576, n_2457);
  not g4678 (n_2458, n2861);
  and g4679 (n2862, n1837, n_2458);
  not g4680 (n_2459, n2862);
  and g4681 (n2863, n1068, n_2459);
  not g4682 (n_2460, n2863);
  and g4683 (n2864, n1072, n_2460);
  not g4684 (n_2461, n2864);
  and g4685 (n2865, n1076, n_2461);
  not g4686 (n_2462, n2865);
  and g4687 (n2866, n1080, n_2462);
  not g4688 (n_2463, n2866);
  and g4689 (n2867, n1084, n_2463);
  not g4690 (n_2464, n2867);
  and g4691 (n2868, n1088, n_2464);
  not g4692 (n_2465, n2868);
  and g4693 (n2869, n1092, n_2465);
  not g4694 (n_2466, n2869);
  and g4695 (n2870, n1096, n_2466);
  not g4696 (n_2467, n2870);
  and g4697 (n2871, n1100, n_2467);
  and g4698 (n2872, \req[19] , n_871);
  not g4699 (n_2468, n2871);
  and g4700 (\grant[19] , n_2468, n2872);
  not g4701 (n_2469, n439);
  and g4702 (n2874, n_2469, n1111);
  not g4703 (n_2470, n2874);
  and g4704 (n2875, n1116, n_2470);
  not g4705 (n_2471, n2875);
  and g4706 (n2876, n1120, n_2471);
  not g4707 (n_2472, n2876);
  and g4708 (n2877, n1124, n_2472);
  not g4709 (n_2473, n2877);
  and g4710 (n2878, n1128, n_2473);
  not g4711 (n_2474, n2878);
  and g4712 (n2879, n1132, n_2474);
  not g4713 (n_2475, n2879);
  and g4714 (n2880, n1136, n_2475);
  not g4715 (n_2476, n2880);
  and g4716 (n2881, n1140, n_2476);
  not g4717 (n_2477, n2881);
  and g4718 (n2882, n1144, n_2477);
  not g4719 (n_2478, n2882);
  and g4720 (n2883, n1148, n_2478);
  not g4721 (n_2479, n2883);
  and g4722 (n2884, n1152, n_2479);
  not g4723 (n_2480, n2884);
  and g4724 (n2885, n1156, n_2480);
  not g4725 (n_2481, n2885);
  and g4726 (n2886, n1160, n_2481);
  not g4727 (n_2482, n2886);
  and g4728 (n2887, n1164, n_2482);
  not g4729 (n_2483, n2887);
  and g4730 (n2888, n1168, n_2483);
  not g4731 (n_2484, n2888);
  and g4732 (n2889, n1172, n_2484);
  not g4733 (n_2485, n2889);
  and g4734 (n2890, n1176, n_2485);
  not g4735 (n_2486, n2890);
  and g4736 (n2891, n1180, n_2486);
  not g4737 (n_2487, n2891);
  and g4738 (n2892, n1184, n_2487);
  not g4739 (n_2488, n2892);
  and g4740 (n2893, n1188, n_2488);
  not g4741 (n_2489, n2893);
  and g4742 (n2894, n1192, n_2489);
  not g4743 (n_2490, n2894);
  and g4744 (n2895, n1196, n_2490);
  not g4745 (n_2491, n2895);
  and g4746 (n2896, n1200, n_2491);
  not g4747 (n_2492, n2896);
  and g4748 (n2897, n1204, n_2492);
  not g4749 (n_2493, n2897);
  and g4750 (n2898, n1208, n_2493);
  not g4751 (n_2494, n2898);
  and g4752 (n2899, n1212, n_2494);
  not g4753 (n_2495, n2899);
  and g4754 (n2900, n1216, n_2495);
  not g4755 (n_2496, n2900);
  and g4756 (n2901, n1220, n_2496);
  not g4757 (n_2497, n2901);
  and g4758 (n2902, n1224, n_2497);
  not g4759 (n_2498, n2902);
  and g4760 (n2903, n1228, n_2498);
  not g4761 (n_2499, n2903);
  and g4762 (n2904, n1232, n_2499);
  not g4763 (n_2500, n2904);
  and g4764 (n2905, n1236, n_2500);
  not g4765 (n_2501, n2905);
  and g4766 (n2906, n1240, n_2501);
  not g4767 (n_2502, n2906);
  and g4768 (n2907, n1244, n_2502);
  not g4769 (n_2503, n2907);
  and g4770 (n2908, n1248, n_2503);
  not g4771 (n_2504, n2908);
  and g4772 (n2909, n1252, n_2504);
  not g4773 (n_2505, n2909);
  and g4774 (n2910, n1256, n_2505);
  not g4775 (n_2506, n2910);
  and g4776 (n2911, n1260, n_2506);
  not g4777 (n_2507, n2911);
  and g4778 (n2912, n1264, n_2507);
  not g4779 (n_2508, n2912);
  and g4780 (n2913, n1268, n_2508);
  not g4781 (n_2509, n2913);
  and g4782 (n2914, n1272, n_2509);
  not g4783 (n_2510, n2914);
  and g4784 (n2915, n1276, n_2510);
  not g4785 (n_2511, n2915);
  and g4786 (n2916, n1280, n_2511);
  not g4787 (n_2512, n2916);
  and g4788 (n2917, n1284, n_2512);
  not g4789 (n_2513, n2917);
  and g4790 (n2918, n1288, n_2513);
  not g4791 (n_2514, n2918);
  and g4792 (n2919, n1292, n_2514);
  not g4793 (n_2515, n2919);
  and g4794 (n2920, n1296, n_2515);
  not g4795 (n_2516, n2920);
  and g4796 (n2921, n1300, n_2516);
  not g4797 (n_2517, n2921);
  and g4798 (n2922, n1304, n_2517);
  not g4799 (n_2518, n2922);
  and g4800 (n2923, n1308, n_2518);
  not g4801 (n_2519, n2923);
  and g4802 (n2924, n1312, n_2519);
  not g4803 (n_2520, n2924);
  and g4804 (n2925, n1316, n_2520);
  not g4805 (n_2521, n2925);
  and g4806 (n2926, n1320, n_2521);
  not g4807 (n_2522, n2926);
  and g4808 (n2927, n1324, n_2522);
  not g4809 (n_2523, n2927);
  and g4810 (n2928, n1328, n_2523);
  not g4811 (n_2524, n2928);
  and g4812 (n2929, n1332, n_2524);
  not g4813 (n_2525, n2929);
  and g4814 (n2930, n1336, n_2525);
  not g4815 (n_2526, n2930);
  and g4816 (n2931, n1340, n_2526);
  not g4817 (n_2527, n2931);
  and g4818 (n2932, n1344, n_2527);
  not g4819 (n_2528, n2932);
  and g4820 (n2933, n1348, n_2528);
  not g4821 (n_2529, n2933);
  and g4822 (n2934, n1352, n_2529);
  not g4823 (n_2530, n2934);
  and g4824 (n2935, n1356, n_2530);
  not g4825 (n_2531, n2935);
  and g4826 (n2936, n1360, n_2531);
  not g4827 (n_2532, n2936);
  and g4828 (n2937, n1364, n_2532);
  not g4829 (n_2533, n2937);
  and g4830 (n2938, n1368, n_2533);
  not g4831 (n_2534, n2938);
  and g4832 (n2939, n1372, n_2534);
  not g4833 (n_2535, n2939);
  and g4834 (n2940, n1376, n_2535);
  not g4835 (n_2536, n2940);
  and g4836 (n2941, n1380, n_2536);
  not g4837 (n_2537, n2941);
  and g4838 (n2942, n1384, n_2537);
  not g4839 (n_2538, n2942);
  and g4840 (n2943, n1388, n_2538);
  not g4841 (n_2539, n2943);
  and g4842 (n2944, n1392, n_2539);
  not g4843 (n_2540, n2944);
  and g4844 (n2945, n1396, n_2540);
  not g4845 (n_2541, n2945);
  and g4846 (n2946, n1663, n_2541);
  not g4847 (n_2542, n2946);
  and g4848 (n2947, n392, n_2542);
  not g4849 (n_2543, n2947);
  and g4850 (n2948, n396, n_2543);
  not g4851 (n_2544, n2948);
  and g4852 (n2949, n400, n_2544);
  not g4853 (n_2545, n2949);
  and g4854 (n2950, n404, n_2545);
  not g4855 (n_2546, n2950);
  and g4856 (n2951, n408, n_2546);
  not g4857 (n_2547, n2951);
  and g4858 (n2952, n412, n_2547);
  not g4859 (n_2548, n2952);
  and g4860 (n2953, n416, n_2548);
  not g4861 (n_2549, n2953);
  and g4862 (n2954, n420, n_2549);
  not g4863 (n_2550, n2954);
  and g4864 (n2955, n424, n_2550);
  not g4865 (n_2551, n2955);
  and g4866 (n2956, n428, n_2551);
  not g4867 (n_2552, n2956);
  and g4868 (n2957, n432, n_2552);
  and g4869 (n2958, \req[20] , n_94);
  not g4870 (n_2553, n2957);
  and g4871 (\grant[20] , n_2553, n2958);
  not g4872 (n_2554, n778);
  and g4873 (n2960, n443, n_2554);
  not g4874 (n_2555, n2960);
  and g4875 (n2961, n448, n_2555);
  not g4876 (n_2556, n2961);
  and g4877 (n2962, n452, n_2556);
  not g4878 (n_2557, n2962);
  and g4879 (n2963, n456, n_2557);
  not g4880 (n_2558, n2963);
  and g4881 (n2964, n460, n_2558);
  not g4882 (n_2559, n2964);
  and g4883 (n2965, n464, n_2559);
  not g4884 (n_2560, n2965);
  and g4885 (n2966, n468, n_2560);
  not g4886 (n_2561, n2966);
  and g4887 (n2967, n472, n_2561);
  not g4888 (n_2562, n2967);
  and g4889 (n2968, n476, n_2562);
  not g4890 (n_2563, n2968);
  and g4891 (n2969, n480, n_2563);
  not g4892 (n_2564, n2969);
  and g4893 (n2970, n484, n_2564);
  not g4894 (n_2565, n2970);
  and g4895 (n2971, n488, n_2565);
  not g4896 (n_2566, n2971);
  and g4897 (n2972, n492, n_2566);
  not g4898 (n_2567, n2972);
  and g4899 (n2973, n496, n_2567);
  not g4900 (n_2568, n2973);
  and g4901 (n2974, n500, n_2568);
  not g4902 (n_2569, n2974);
  and g4903 (n2975, n504, n_2569);
  not g4904 (n_2570, n2975);
  and g4905 (n2976, n508, n_2570);
  not g4906 (n_2571, n2976);
  and g4907 (n2977, n512, n_2571);
  not g4908 (n_2572, n2977);
  and g4909 (n2978, n516, n_2572);
  not g4910 (n_2573, n2978);
  and g4911 (n2979, n520, n_2573);
  not g4912 (n_2574, n2979);
  and g4913 (n2980, n524, n_2574);
  not g4914 (n_2575, n2980);
  and g4915 (n2981, n528, n_2575);
  not g4916 (n_2576, n2981);
  and g4917 (n2982, n532, n_2576);
  not g4918 (n_2577, n2982);
  and g4919 (n2983, n536, n_2577);
  not g4920 (n_2578, n2983);
  and g4921 (n2984, n540, n_2578);
  not g4922 (n_2579, n2984);
  and g4923 (n2985, n544, n_2579);
  not g4924 (n_2580, n2985);
  and g4925 (n2986, n548, n_2580);
  not g4926 (n_2581, n2986);
  and g4927 (n2987, n552, n_2581);
  not g4928 (n_2582, n2987);
  and g4929 (n2988, n556, n_2582);
  not g4930 (n_2583, n2988);
  and g4931 (n2989, n560, n_2583);
  not g4932 (n_2584, n2989);
  and g4933 (n2990, n564, n_2584);
  not g4934 (n_2585, n2990);
  and g4935 (n2991, n568, n_2585);
  not g4936 (n_2586, n2991);
  and g4937 (n2992, n572, n_2586);
  not g4938 (n_2587, n2992);
  and g4939 (n2993, n576, n_2587);
  not g4940 (n_2588, n2993);
  and g4941 (n2994, n580, n_2588);
  not g4942 (n_2589, n2994);
  and g4943 (n2995, n584, n_2589);
  not g4944 (n_2590, n2995);
  and g4945 (n2996, n588, n_2590);
  not g4946 (n_2591, n2996);
  and g4947 (n2997, n592, n_2591);
  not g4948 (n_2592, n2997);
  and g4949 (n2998, n596, n_2592);
  not g4950 (n_2593, n2998);
  and g4951 (n2999, n600, n_2593);
  not g4952 (n_2594, n2999);
  and g4953 (n3000, n604, n_2594);
  not g4954 (n_2595, n3000);
  and g4955 (n3001, n608, n_2595);
  not g4956 (n_2596, n3001);
  and g4957 (n3002, n612, n_2596);
  not g4958 (n_2597, n3002);
  and g4959 (n3003, n616, n_2597);
  not g4960 (n_2598, n3003);
  and g4961 (n3004, n620, n_2598);
  not g4962 (n_2599, n3004);
  and g4963 (n3005, n624, n_2599);
  not g4964 (n_2600, n3005);
  and g4965 (n3006, n628, n_2600);
  not g4966 (n_2601, n3006);
  and g4967 (n3007, n632, n_2601);
  not g4968 (n_2602, n3007);
  and g4969 (n3008, n636, n_2602);
  not g4970 (n_2603, n3008);
  and g4971 (n3009, n640, n_2603);
  not g4972 (n_2604, n3009);
  and g4973 (n3010, n644, n_2604);
  not g4974 (n_2605, n3010);
  and g4975 (n3011, n648, n_2605);
  not g4976 (n_2606, n3011);
  and g4977 (n3012, n652, n_2606);
  not g4978 (n_2607, n3012);
  and g4979 (n3013, n656, n_2607);
  not g4980 (n_2608, n3013);
  and g4981 (n3014, n660, n_2608);
  not g4982 (n_2609, n3014);
  and g4983 (n3015, n664, n_2609);
  not g4984 (n_2610, n3015);
  and g4985 (n3016, n668, n_2610);
  not g4986 (n_2611, n3016);
  and g4987 (n3017, n672, n_2611);
  not g4988 (n_2612, n3017);
  and g4989 (n3018, n676, n_2612);
  not g4990 (n_2613, n3018);
  and g4991 (n3019, n680, n_2613);
  not g4992 (n_2614, n3019);
  and g4993 (n3020, n684, n_2614);
  not g4994 (n_2615, n3020);
  and g4995 (n3021, n688, n_2615);
  not g4996 (n_2616, n3021);
  and g4997 (n3022, n692, n_2616);
  not g4998 (n_2617, n3022);
  and g4999 (n3023, n696, n_2617);
  not g5000 (n_2618, n3023);
  and g5001 (n3024, n700, n_2618);
  not g5002 (n_2619, n3024);
  and g5003 (n3025, n704, n_2619);
  not g5004 (n_2620, n3025);
  and g5005 (n3026, n708, n_2620);
  not g5006 (n_2621, n3026);
  and g5007 (n3027, n712, n_2621);
  not g5008 (n_2622, n3027);
  and g5009 (n3028, n716, n_2622);
  not g5010 (n_2623, n3028);
  and g5011 (n3029, n720, n_2623);
  not g5012 (n_2624, n3029);
  and g5013 (n3030, n1484, n_2624);
  not g5014 (n_2625, n3030);
  and g5015 (n3031, n1486, n_2625);
  not g5016 (n_2626, n3031);
  and g5017 (n3032, n1750, n_2626);
  not g5018 (n_2627, n3032);
  and g5019 (n3033, n731, n_2627);
  not g5020 (n_2628, n3033);
  and g5021 (n3034, n735, n_2628);
  not g5022 (n_2629, n3034);
  and g5023 (n3035, n739, n_2629);
  not g5024 (n_2630, n3035);
  and g5025 (n3036, n743, n_2630);
  not g5026 (n_2631, n3036);
  and g5027 (n3037, n747, n_2631);
  not g5028 (n_2632, n3037);
  and g5029 (n3038, n751, n_2632);
  not g5030 (n_2633, n3038);
  and g5031 (n3039, n755, n_2633);
  not g5032 (n_2634, n3039);
  and g5033 (n3040, n759, n_2634);
  not g5034 (n_2635, n3040);
  and g5035 (n3041, n763, n_2635);
  not g5036 (n_2636, n3041);
  and g5037 (n3042, n767, n_2636);
  not g5038 (n_2637, n3042);
  and g5039 (n3043, n771, n_2637);
  and g5040 (n3044, \req[21] , n_635);
  not g5041 (n_2638, n3043);
  and g5042 (\grant[21] , n_2638, n3044);
  not g5043 (n_2639, n1115);
  and g5044 (n3046, n782, n_2639);
  not g5045 (n_2640, n3046);
  and g5046 (n3047, n787, n_2640);
  not g5047 (n_2641, n3047);
  and g5048 (n3048, n791, n_2641);
  not g5049 (n_2642, n3048);
  and g5050 (n3049, n795, n_2642);
  not g5051 (n_2643, n3049);
  and g5052 (n3050, n799, n_2643);
  not g5053 (n_2644, n3050);
  and g5054 (n3051, n803, n_2644);
  not g5055 (n_2645, n3051);
  and g5056 (n3052, n807, n_2645);
  not g5057 (n_2646, n3052);
  and g5058 (n3053, n811, n_2646);
  not g5059 (n_2647, n3053);
  and g5060 (n3054, n815, n_2647);
  not g5061 (n_2648, n3054);
  and g5062 (n3055, n819, n_2648);
  not g5063 (n_2649, n3055);
  and g5064 (n3056, n823, n_2649);
  not g5065 (n_2650, n3056);
  and g5066 (n3057, n827, n_2650);
  not g5067 (n_2651, n3057);
  and g5068 (n3058, n831, n_2651);
  not g5069 (n_2652, n3058);
  and g5070 (n3059, n835, n_2652);
  not g5071 (n_2653, n3059);
  and g5072 (n3060, n839, n_2653);
  not g5073 (n_2654, n3060);
  and g5074 (n3061, n843, n_2654);
  not g5075 (n_2655, n3061);
  and g5076 (n3062, n847, n_2655);
  not g5077 (n_2656, n3062);
  and g5078 (n3063, n851, n_2656);
  not g5079 (n_2657, n3063);
  and g5080 (n3064, n855, n_2657);
  not g5081 (n_2658, n3064);
  and g5082 (n3065, n859, n_2658);
  not g5083 (n_2659, n3065);
  and g5084 (n3066, n863, n_2659);
  not g5085 (n_2660, n3066);
  and g5086 (n3067, n867, n_2660);
  not g5087 (n_2661, n3067);
  and g5088 (n3068, n871, n_2661);
  not g5089 (n_2662, n3068);
  and g5090 (n3069, n875, n_2662);
  not g5091 (n_2663, n3069);
  and g5092 (n3070, n879, n_2663);
  not g5093 (n_2664, n3070);
  and g5094 (n3071, n883, n_2664);
  not g5095 (n_2665, n3071);
  and g5096 (n3072, n887, n_2665);
  not g5097 (n_2666, n3072);
  and g5098 (n3073, n891, n_2666);
  not g5099 (n_2667, n3073);
  and g5100 (n3074, n895, n_2667);
  not g5101 (n_2668, n3074);
  and g5102 (n3075, n899, n_2668);
  not g5103 (n_2669, n3075);
  and g5104 (n3076, n903, n_2669);
  not g5105 (n_2670, n3076);
  and g5106 (n3077, n907, n_2670);
  not g5107 (n_2671, n3077);
  and g5108 (n3078, n911, n_2671);
  not g5109 (n_2672, n3078);
  and g5110 (n3079, n915, n_2672);
  not g5111 (n_2673, n3079);
  and g5112 (n3080, n919, n_2673);
  not g5113 (n_2674, n3080);
  and g5114 (n3081, n923, n_2674);
  not g5115 (n_2675, n3081);
  and g5116 (n3082, n927, n_2675);
  not g5117 (n_2676, n3082);
  and g5118 (n3083, n931, n_2676);
  not g5119 (n_2677, n3083);
  and g5120 (n3084, n935, n_2677);
  not g5121 (n_2678, n3084);
  and g5122 (n3085, n939, n_2678);
  not g5123 (n_2679, n3085);
  and g5124 (n3086, n943, n_2679);
  not g5125 (n_2680, n3086);
  and g5126 (n3087, n947, n_2680);
  not g5127 (n_2681, n3087);
  and g5128 (n3088, n951, n_2681);
  not g5129 (n_2682, n3088);
  and g5130 (n3089, n955, n_2682);
  not g5131 (n_2683, n3089);
  and g5132 (n3090, n959, n_2683);
  not g5133 (n_2684, n3090);
  and g5134 (n3091, n963, n_2684);
  not g5135 (n_2685, n3091);
  and g5136 (n3092, n967, n_2685);
  not g5137 (n_2686, n3092);
  and g5138 (n3093, n971, n_2686);
  not g5139 (n_2687, n3093);
  and g5140 (n3094, n975, n_2687);
  not g5141 (n_2688, n3094);
  and g5142 (n3095, n979, n_2688);
  not g5143 (n_2689, n3095);
  and g5144 (n3096, n983, n_2689);
  not g5145 (n_2690, n3096);
  and g5146 (n3097, n987, n_2690);
  not g5147 (n_2691, n3097);
  and g5148 (n3098, n991, n_2691);
  not g5149 (n_2692, n3098);
  and g5150 (n3099, n995, n_2692);
  not g5151 (n_2693, n3099);
  and g5152 (n3100, n999, n_2693);
  not g5153 (n_2694, n3100);
  and g5154 (n3101, n1003, n_2694);
  not g5155 (n_2695, n3101);
  and g5156 (n3102, n1007, n_2695);
  not g5157 (n_2696, n3102);
  and g5158 (n3103, n1011, n_2696);
  not g5159 (n_2697, n3103);
  and g5160 (n3104, n1015, n_2697);
  not g5161 (n_2698, n3104);
  and g5162 (n3105, n1019, n_2698);
  not g5163 (n_2699, n3105);
  and g5164 (n3106, n1023, n_2699);
  not g5165 (n_2700, n3106);
  and g5166 (n3107, n1027, n_2700);
  not g5167 (n_2701, n3107);
  and g5168 (n3108, n1031, n_2701);
  not g5169 (n_2702, n3108);
  and g5170 (n3109, n1035, n_2702);
  not g5171 (n_2703, n3109);
  and g5172 (n3110, n1039, n_2703);
  not g5173 (n_2704, n3110);
  and g5174 (n3111, n1043, n_2704);
  not g5175 (n_2705, n3111);
  and g5176 (n3112, n1047, n_2705);
  not g5177 (n_2706, n3112);
  and g5178 (n3113, n1051, n_2706);
  not g5179 (n_2707, n3113);
  and g5180 (n3114, n1055, n_2707);
  not g5181 (n_2708, n3114);
  and g5182 (n3115, n1059, n_2708);
  not g5183 (n_2709, n3115);
  and g5184 (n3116, n1574, n_2709);
  not g5185 (n_2710, n3116);
  and g5186 (n3117, n1576, n_2710);
  not g5187 (n_2711, n3117);
  and g5188 (n3118, n1837, n_2711);
  not g5189 (n_2712, n3118);
  and g5190 (n3119, n1068, n_2712);
  not g5191 (n_2713, n3119);
  and g5192 (n3120, n1072, n_2713);
  not g5193 (n_2714, n3120);
  and g5194 (n3121, n1076, n_2714);
  not g5195 (n_2715, n3121);
  and g5196 (n3122, n1080, n_2715);
  not g5197 (n_2716, n3122);
  and g5198 (n3123, n1084, n_2716);
  not g5199 (n_2717, n3123);
  and g5200 (n3124, n1088, n_2717);
  not g5201 (n_2718, n3124);
  and g5202 (n3125, n1092, n_2718);
  not g5203 (n_2719, n3125);
  and g5204 (n3126, n1096, n_2719);
  not g5205 (n_2720, n3126);
  and g5206 (n3127, n1100, n_2720);
  not g5207 (n_2721, n3127);
  and g5208 (n3128, n1104, n_2721);
  not g5209 (n_2722, n3128);
  and g5210 (n3129, n1108, n_2722);
  and g5211 (n3130, \req[22] , n_875);
  not g5212 (n_2723, n3129);
  and g5213 (\grant[22] , n_2723, n3130);
  not g5214 (n_2724, n447);
  and g5215 (n3132, n_2724, n1119);
  not g5216 (n_2725, n3132);
  and g5217 (n3133, n1124, n_2725);
  not g5218 (n_2726, n3133);
  and g5219 (n3134, n1128, n_2726);
  not g5220 (n_2727, n3134);
  and g5221 (n3135, n1132, n_2727);
  not g5222 (n_2728, n3135);
  and g5223 (n3136, n1136, n_2728);
  not g5224 (n_2729, n3136);
  and g5225 (n3137, n1140, n_2729);
  not g5226 (n_2730, n3137);
  and g5227 (n3138, n1144, n_2730);
  not g5228 (n_2731, n3138);
  and g5229 (n3139, n1148, n_2731);
  not g5230 (n_2732, n3139);
  and g5231 (n3140, n1152, n_2732);
  not g5232 (n_2733, n3140);
  and g5233 (n3141, n1156, n_2733);
  not g5234 (n_2734, n3141);
  and g5235 (n3142, n1160, n_2734);
  not g5236 (n_2735, n3142);
  and g5237 (n3143, n1164, n_2735);
  not g5238 (n_2736, n3143);
  and g5239 (n3144, n1168, n_2736);
  not g5240 (n_2737, n3144);
  and g5241 (n3145, n1172, n_2737);
  not g5242 (n_2738, n3145);
  and g5243 (n3146, n1176, n_2738);
  not g5244 (n_2739, n3146);
  and g5245 (n3147, n1180, n_2739);
  not g5246 (n_2740, n3147);
  and g5247 (n3148, n1184, n_2740);
  not g5248 (n_2741, n3148);
  and g5249 (n3149, n1188, n_2741);
  not g5250 (n_2742, n3149);
  and g5251 (n3150, n1192, n_2742);
  not g5252 (n_2743, n3150);
  and g5253 (n3151, n1196, n_2743);
  not g5254 (n_2744, n3151);
  and g5255 (n3152, n1200, n_2744);
  not g5256 (n_2745, n3152);
  and g5257 (n3153, n1204, n_2745);
  not g5258 (n_2746, n3153);
  and g5259 (n3154, n1208, n_2746);
  not g5260 (n_2747, n3154);
  and g5261 (n3155, n1212, n_2747);
  not g5262 (n_2748, n3155);
  and g5263 (n3156, n1216, n_2748);
  not g5264 (n_2749, n3156);
  and g5265 (n3157, n1220, n_2749);
  not g5266 (n_2750, n3157);
  and g5267 (n3158, n1224, n_2750);
  not g5268 (n_2751, n3158);
  and g5269 (n3159, n1228, n_2751);
  not g5270 (n_2752, n3159);
  and g5271 (n3160, n1232, n_2752);
  not g5272 (n_2753, n3160);
  and g5273 (n3161, n1236, n_2753);
  not g5274 (n_2754, n3161);
  and g5275 (n3162, n1240, n_2754);
  not g5276 (n_2755, n3162);
  and g5277 (n3163, n1244, n_2755);
  not g5278 (n_2756, n3163);
  and g5279 (n3164, n1248, n_2756);
  not g5280 (n_2757, n3164);
  and g5281 (n3165, n1252, n_2757);
  not g5282 (n_2758, n3165);
  and g5283 (n3166, n1256, n_2758);
  not g5284 (n_2759, n3166);
  and g5285 (n3167, n1260, n_2759);
  not g5286 (n_2760, n3167);
  and g5287 (n3168, n1264, n_2760);
  not g5288 (n_2761, n3168);
  and g5289 (n3169, n1268, n_2761);
  not g5290 (n_2762, n3169);
  and g5291 (n3170, n1272, n_2762);
  not g5292 (n_2763, n3170);
  and g5293 (n3171, n1276, n_2763);
  not g5294 (n_2764, n3171);
  and g5295 (n3172, n1280, n_2764);
  not g5296 (n_2765, n3172);
  and g5297 (n3173, n1284, n_2765);
  not g5298 (n_2766, n3173);
  and g5299 (n3174, n1288, n_2766);
  not g5300 (n_2767, n3174);
  and g5301 (n3175, n1292, n_2767);
  not g5302 (n_2768, n3175);
  and g5303 (n3176, n1296, n_2768);
  not g5304 (n_2769, n3176);
  and g5305 (n3177, n1300, n_2769);
  not g5306 (n_2770, n3177);
  and g5307 (n3178, n1304, n_2770);
  not g5308 (n_2771, n3178);
  and g5309 (n3179, n1308, n_2771);
  not g5310 (n_2772, n3179);
  and g5311 (n3180, n1312, n_2772);
  not g5312 (n_2773, n3180);
  and g5313 (n3181, n1316, n_2773);
  not g5314 (n_2774, n3181);
  and g5315 (n3182, n1320, n_2774);
  not g5316 (n_2775, n3182);
  and g5317 (n3183, n1324, n_2775);
  not g5318 (n_2776, n3183);
  and g5319 (n3184, n1328, n_2776);
  not g5320 (n_2777, n3184);
  and g5321 (n3185, n1332, n_2777);
  not g5322 (n_2778, n3185);
  and g5323 (n3186, n1336, n_2778);
  not g5324 (n_2779, n3186);
  and g5325 (n3187, n1340, n_2779);
  not g5326 (n_2780, n3187);
  and g5327 (n3188, n1344, n_2780);
  not g5328 (n_2781, n3188);
  and g5329 (n3189, n1348, n_2781);
  not g5330 (n_2782, n3189);
  and g5331 (n3190, n1352, n_2782);
  not g5332 (n_2783, n3190);
  and g5333 (n3191, n1356, n_2783);
  not g5334 (n_2784, n3191);
  and g5335 (n3192, n1360, n_2784);
  not g5336 (n_2785, n3192);
  and g5337 (n3193, n1364, n_2785);
  not g5338 (n_2786, n3193);
  and g5339 (n3194, n1368, n_2786);
  not g5340 (n_2787, n3194);
  and g5341 (n3195, n1372, n_2787);
  not g5342 (n_2788, n3195);
  and g5343 (n3196, n1376, n_2788);
  not g5344 (n_2789, n3196);
  and g5345 (n3197, n1380, n_2789);
  not g5346 (n_2790, n3197);
  and g5347 (n3198, n1384, n_2790);
  not g5348 (n_2791, n3198);
  and g5349 (n3199, n1388, n_2791);
  not g5350 (n_2792, n3199);
  and g5351 (n3200, n1392, n_2792);
  not g5352 (n_2793, n3200);
  and g5353 (n3201, n1396, n_2793);
  not g5354 (n_2794, n3201);
  and g5355 (n3202, n1663, n_2794);
  not g5356 (n_2795, n3202);
  and g5357 (n3203, n392, n_2795);
  not g5358 (n_2796, n3203);
  and g5359 (n3204, n396, n_2796);
  not g5360 (n_2797, n3204);
  and g5361 (n3205, n400, n_2797);
  not g5362 (n_2798, n3205);
  and g5363 (n3206, n404, n_2798);
  not g5364 (n_2799, n3206);
  and g5365 (n3207, n408, n_2799);
  not g5366 (n_2800, n3207);
  and g5367 (n3208, n412, n_2800);
  not g5368 (n_2801, n3208);
  and g5369 (n3209, n416, n_2801);
  not g5370 (n_2802, n3209);
  and g5371 (n3210, n420, n_2802);
  not g5372 (n_2803, n3210);
  and g5373 (n3211, n424, n_2803);
  not g5374 (n_2804, n3211);
  and g5375 (n3212, n428, n_2804);
  not g5376 (n_2805, n3212);
  and g5377 (n3213, n432, n_2805);
  not g5378 (n_2806, n3213);
  and g5379 (n3214, n436, n_2806);
  not g5380 (n_2807, n3214);
  and g5381 (n3215, n440, n_2807);
  and g5382 (n3216, \req[23] , n_108);
  not g5383 (n_2808, n3215);
  and g5384 (\grant[23] , n_2808, n3216);
  not g5385 (n_2809, n786);
  and g5386 (n3218, n451, n_2809);
  not g5387 (n_2810, n3218);
  and g5388 (n3219, n456, n_2810);
  not g5389 (n_2811, n3219);
  and g5390 (n3220, n460, n_2811);
  not g5391 (n_2812, n3220);
  and g5392 (n3221, n464, n_2812);
  not g5393 (n_2813, n3221);
  and g5394 (n3222, n468, n_2813);
  not g5395 (n_2814, n3222);
  and g5396 (n3223, n472, n_2814);
  not g5397 (n_2815, n3223);
  and g5398 (n3224, n476, n_2815);
  not g5399 (n_2816, n3224);
  and g5400 (n3225, n480, n_2816);
  not g5401 (n_2817, n3225);
  and g5402 (n3226, n484, n_2817);
  not g5403 (n_2818, n3226);
  and g5404 (n3227, n488, n_2818);
  not g5405 (n_2819, n3227);
  and g5406 (n3228, n492, n_2819);
  not g5407 (n_2820, n3228);
  and g5408 (n3229, n496, n_2820);
  not g5409 (n_2821, n3229);
  and g5410 (n3230, n500, n_2821);
  not g5411 (n_2822, n3230);
  and g5412 (n3231, n504, n_2822);
  not g5413 (n_2823, n3231);
  and g5414 (n3232, n508, n_2823);
  not g5415 (n_2824, n3232);
  and g5416 (n3233, n512, n_2824);
  not g5417 (n_2825, n3233);
  and g5418 (n3234, n516, n_2825);
  not g5419 (n_2826, n3234);
  and g5420 (n3235, n520, n_2826);
  not g5421 (n_2827, n3235);
  and g5422 (n3236, n524, n_2827);
  not g5423 (n_2828, n3236);
  and g5424 (n3237, n528, n_2828);
  not g5425 (n_2829, n3237);
  and g5426 (n3238, n532, n_2829);
  not g5427 (n_2830, n3238);
  and g5428 (n3239, n536, n_2830);
  not g5429 (n_2831, n3239);
  and g5430 (n3240, n540, n_2831);
  not g5431 (n_2832, n3240);
  and g5432 (n3241, n544, n_2832);
  not g5433 (n_2833, n3241);
  and g5434 (n3242, n548, n_2833);
  not g5435 (n_2834, n3242);
  and g5436 (n3243, n552, n_2834);
  not g5437 (n_2835, n3243);
  and g5438 (n3244, n556, n_2835);
  not g5439 (n_2836, n3244);
  and g5440 (n3245, n560, n_2836);
  not g5441 (n_2837, n3245);
  and g5442 (n3246, n564, n_2837);
  not g5443 (n_2838, n3246);
  and g5444 (n3247, n568, n_2838);
  not g5445 (n_2839, n3247);
  and g5446 (n3248, n572, n_2839);
  not g5447 (n_2840, n3248);
  and g5448 (n3249, n576, n_2840);
  not g5449 (n_2841, n3249);
  and g5450 (n3250, n580, n_2841);
  not g5451 (n_2842, n3250);
  and g5452 (n3251, n584, n_2842);
  not g5453 (n_2843, n3251);
  and g5454 (n3252, n588, n_2843);
  not g5455 (n_2844, n3252);
  and g5456 (n3253, n592, n_2844);
  not g5457 (n_2845, n3253);
  and g5458 (n3254, n596, n_2845);
  not g5459 (n_2846, n3254);
  and g5460 (n3255, n600, n_2846);
  not g5461 (n_2847, n3255);
  and g5462 (n3256, n604, n_2847);
  not g5463 (n_2848, n3256);
  and g5464 (n3257, n608, n_2848);
  not g5465 (n_2849, n3257);
  and g5466 (n3258, n612, n_2849);
  not g5467 (n_2850, n3258);
  and g5468 (n3259, n616, n_2850);
  not g5469 (n_2851, n3259);
  and g5470 (n3260, n620, n_2851);
  not g5471 (n_2852, n3260);
  and g5472 (n3261, n624, n_2852);
  not g5473 (n_2853, n3261);
  and g5474 (n3262, n628, n_2853);
  not g5475 (n_2854, n3262);
  and g5476 (n3263, n632, n_2854);
  not g5477 (n_2855, n3263);
  and g5478 (n3264, n636, n_2855);
  not g5479 (n_2856, n3264);
  and g5480 (n3265, n640, n_2856);
  not g5481 (n_2857, n3265);
  and g5482 (n3266, n644, n_2857);
  not g5483 (n_2858, n3266);
  and g5484 (n3267, n648, n_2858);
  not g5485 (n_2859, n3267);
  and g5486 (n3268, n652, n_2859);
  not g5487 (n_2860, n3268);
  and g5488 (n3269, n656, n_2860);
  not g5489 (n_2861, n3269);
  and g5490 (n3270, n660, n_2861);
  not g5491 (n_2862, n3270);
  and g5492 (n3271, n664, n_2862);
  not g5493 (n_2863, n3271);
  and g5494 (n3272, n668, n_2863);
  not g5495 (n_2864, n3272);
  and g5496 (n3273, n672, n_2864);
  not g5497 (n_2865, n3273);
  and g5498 (n3274, n676, n_2865);
  not g5499 (n_2866, n3274);
  and g5500 (n3275, n680, n_2866);
  not g5501 (n_2867, n3275);
  and g5502 (n3276, n684, n_2867);
  not g5503 (n_2868, n3276);
  and g5504 (n3277, n688, n_2868);
  not g5505 (n_2869, n3277);
  and g5506 (n3278, n692, n_2869);
  not g5507 (n_2870, n3278);
  and g5508 (n3279, n696, n_2870);
  not g5509 (n_2871, n3279);
  and g5510 (n3280, n700, n_2871);
  not g5511 (n_2872, n3280);
  and g5512 (n3281, n704, n_2872);
  not g5513 (n_2873, n3281);
  and g5514 (n3282, n708, n_2873);
  not g5515 (n_2874, n3282);
  and g5516 (n3283, n712, n_2874);
  not g5517 (n_2875, n3283);
  and g5518 (n3284, n716, n_2875);
  not g5519 (n_2876, n3284);
  and g5520 (n3285, n720, n_2876);
  not g5521 (n_2877, n3285);
  and g5522 (n3286, n1484, n_2877);
  not g5523 (n_2878, n3286);
  and g5524 (n3287, n1486, n_2878);
  not g5525 (n_2879, n3287);
  and g5526 (n3288, n1750, n_2879);
  not g5527 (n_2880, n3288);
  and g5528 (n3289, n731, n_2880);
  not g5529 (n_2881, n3289);
  and g5530 (n3290, n735, n_2881);
  not g5531 (n_2882, n3290);
  and g5532 (n3291, n739, n_2882);
  not g5533 (n_2883, n3291);
  and g5534 (n3292, n743, n_2883);
  not g5535 (n_2884, n3292);
  and g5536 (n3293, n747, n_2884);
  not g5537 (n_2885, n3293);
  and g5538 (n3294, n751, n_2885);
  not g5539 (n_2886, n3294);
  and g5540 (n3295, n755, n_2886);
  not g5541 (n_2887, n3295);
  and g5542 (n3296, n759, n_2887);
  not g5543 (n_2888, n3296);
  and g5544 (n3297, n763, n_2888);
  not g5545 (n_2889, n3297);
  and g5546 (n3298, n767, n_2889);
  not g5547 (n_2890, n3298);
  and g5548 (n3299, n771, n_2890);
  not g5549 (n_2891, n3299);
  and g5550 (n3300, n775, n_2891);
  not g5551 (n_2892, n3300);
  and g5552 (n3301, n779, n_2892);
  and g5553 (n3302, \req[24] , n_641);
  not g5554 (n_2893, n3301);
  and g5555 (\grant[24] , n_2893, n3302);
  not g5556 (n_2894, n1123);
  and g5557 (n3304, n790, n_2894);
  not g5558 (n_2895, n3304);
  and g5559 (n3305, n795, n_2895);
  not g5560 (n_2896, n3305);
  and g5561 (n3306, n799, n_2896);
  not g5562 (n_2897, n3306);
  and g5563 (n3307, n803, n_2897);
  not g5564 (n_2898, n3307);
  and g5565 (n3308, n807, n_2898);
  not g5566 (n_2899, n3308);
  and g5567 (n3309, n811, n_2899);
  not g5568 (n_2900, n3309);
  and g5569 (n3310, n815, n_2900);
  not g5570 (n_2901, n3310);
  and g5571 (n3311, n819, n_2901);
  not g5572 (n_2902, n3311);
  and g5573 (n3312, n823, n_2902);
  not g5574 (n_2903, n3312);
  and g5575 (n3313, n827, n_2903);
  not g5576 (n_2904, n3313);
  and g5577 (n3314, n831, n_2904);
  not g5578 (n_2905, n3314);
  and g5579 (n3315, n835, n_2905);
  not g5580 (n_2906, n3315);
  and g5581 (n3316, n839, n_2906);
  not g5582 (n_2907, n3316);
  and g5583 (n3317, n843, n_2907);
  not g5584 (n_2908, n3317);
  and g5585 (n3318, n847, n_2908);
  not g5586 (n_2909, n3318);
  and g5587 (n3319, n851, n_2909);
  not g5588 (n_2910, n3319);
  and g5589 (n3320, n855, n_2910);
  not g5590 (n_2911, n3320);
  and g5591 (n3321, n859, n_2911);
  not g5592 (n_2912, n3321);
  and g5593 (n3322, n863, n_2912);
  not g5594 (n_2913, n3322);
  and g5595 (n3323, n867, n_2913);
  not g5596 (n_2914, n3323);
  and g5597 (n3324, n871, n_2914);
  not g5598 (n_2915, n3324);
  and g5599 (n3325, n875, n_2915);
  not g5600 (n_2916, n3325);
  and g5601 (n3326, n879, n_2916);
  not g5602 (n_2917, n3326);
  and g5603 (n3327, n883, n_2917);
  not g5604 (n_2918, n3327);
  and g5605 (n3328, n887, n_2918);
  not g5606 (n_2919, n3328);
  and g5607 (n3329, n891, n_2919);
  not g5608 (n_2920, n3329);
  and g5609 (n3330, n895, n_2920);
  not g5610 (n_2921, n3330);
  and g5611 (n3331, n899, n_2921);
  not g5612 (n_2922, n3331);
  and g5613 (n3332, n903, n_2922);
  not g5614 (n_2923, n3332);
  and g5615 (n3333, n907, n_2923);
  not g5616 (n_2924, n3333);
  and g5617 (n3334, n911, n_2924);
  not g5618 (n_2925, n3334);
  and g5619 (n3335, n915, n_2925);
  not g5620 (n_2926, n3335);
  and g5621 (n3336, n919, n_2926);
  not g5622 (n_2927, n3336);
  and g5623 (n3337, n923, n_2927);
  not g5624 (n_2928, n3337);
  and g5625 (n3338, n927, n_2928);
  not g5626 (n_2929, n3338);
  and g5627 (n3339, n931, n_2929);
  not g5628 (n_2930, n3339);
  and g5629 (n3340, n935, n_2930);
  not g5630 (n_2931, n3340);
  and g5631 (n3341, n939, n_2931);
  not g5632 (n_2932, n3341);
  and g5633 (n3342, n943, n_2932);
  not g5634 (n_2933, n3342);
  and g5635 (n3343, n947, n_2933);
  not g5636 (n_2934, n3343);
  and g5637 (n3344, n951, n_2934);
  not g5638 (n_2935, n3344);
  and g5639 (n3345, n955, n_2935);
  not g5640 (n_2936, n3345);
  and g5641 (n3346, n959, n_2936);
  not g5642 (n_2937, n3346);
  and g5643 (n3347, n963, n_2937);
  not g5644 (n_2938, n3347);
  and g5645 (n3348, n967, n_2938);
  not g5646 (n_2939, n3348);
  and g5647 (n3349, n971, n_2939);
  not g5648 (n_2940, n3349);
  and g5649 (n3350, n975, n_2940);
  not g5650 (n_2941, n3350);
  and g5651 (n3351, n979, n_2941);
  not g5652 (n_2942, n3351);
  and g5653 (n3352, n983, n_2942);
  not g5654 (n_2943, n3352);
  and g5655 (n3353, n987, n_2943);
  not g5656 (n_2944, n3353);
  and g5657 (n3354, n991, n_2944);
  not g5658 (n_2945, n3354);
  and g5659 (n3355, n995, n_2945);
  not g5660 (n_2946, n3355);
  and g5661 (n3356, n999, n_2946);
  not g5662 (n_2947, n3356);
  and g5663 (n3357, n1003, n_2947);
  not g5664 (n_2948, n3357);
  and g5665 (n3358, n1007, n_2948);
  not g5666 (n_2949, n3358);
  and g5667 (n3359, n1011, n_2949);
  not g5668 (n_2950, n3359);
  and g5669 (n3360, n1015, n_2950);
  not g5670 (n_2951, n3360);
  and g5671 (n3361, n1019, n_2951);
  not g5672 (n_2952, n3361);
  and g5673 (n3362, n1023, n_2952);
  not g5674 (n_2953, n3362);
  and g5675 (n3363, n1027, n_2953);
  not g5676 (n_2954, n3363);
  and g5677 (n3364, n1031, n_2954);
  not g5678 (n_2955, n3364);
  and g5679 (n3365, n1035, n_2955);
  not g5680 (n_2956, n3365);
  and g5681 (n3366, n1039, n_2956);
  not g5682 (n_2957, n3366);
  and g5683 (n3367, n1043, n_2957);
  not g5684 (n_2958, n3367);
  and g5685 (n3368, n1047, n_2958);
  not g5686 (n_2959, n3368);
  and g5687 (n3369, n1051, n_2959);
  not g5688 (n_2960, n3369);
  and g5689 (n3370, n1055, n_2960);
  not g5690 (n_2961, n3370);
  and g5691 (n3371, n1059, n_2961);
  not g5692 (n_2962, n3371);
  and g5693 (n3372, n1574, n_2962);
  not g5694 (n_2963, n3372);
  and g5695 (n3373, n1576, n_2963);
  not g5696 (n_2964, n3373);
  and g5697 (n3374, n1837, n_2964);
  not g5698 (n_2965, n3374);
  and g5699 (n3375, n1068, n_2965);
  not g5700 (n_2966, n3375);
  and g5701 (n3376, n1072, n_2966);
  not g5702 (n_2967, n3376);
  and g5703 (n3377, n1076, n_2967);
  not g5704 (n_2968, n3377);
  and g5705 (n3378, n1080, n_2968);
  not g5706 (n_2969, n3378);
  and g5707 (n3379, n1084, n_2969);
  not g5708 (n_2970, n3379);
  and g5709 (n3380, n1088, n_2970);
  not g5710 (n_2971, n3380);
  and g5711 (n3381, n1092, n_2971);
  not g5712 (n_2972, n3381);
  and g5713 (n3382, n1096, n_2972);
  not g5714 (n_2973, n3382);
  and g5715 (n3383, n1100, n_2973);
  not g5716 (n_2974, n3383);
  and g5717 (n3384, n1104, n_2974);
  not g5718 (n_2975, n3384);
  and g5719 (n3385, n1108, n_2975);
  not g5720 (n_2976, n3385);
  and g5721 (n3386, n1112, n_2976);
  not g5722 (n_2977, n3386);
  and g5723 (n3387, n1116, n_2977);
  and g5724 (n3388, \req[25] , n_879);
  not g5725 (n_2978, n3387);
  and g5726 (\grant[25] , n_2978, n3388);
  not g5727 (n_2979, n455);
  and g5728 (n3390, n_2979, n1127);
  not g5729 (n_2980, n3390);
  and g5730 (n3391, n1132, n_2980);
  not g5731 (n_2981, n3391);
  and g5732 (n3392, n1136, n_2981);
  not g5733 (n_2982, n3392);
  and g5734 (n3393, n1140, n_2982);
  not g5735 (n_2983, n3393);
  and g5736 (n3394, n1144, n_2983);
  not g5737 (n_2984, n3394);
  and g5738 (n3395, n1148, n_2984);
  not g5739 (n_2985, n3395);
  and g5740 (n3396, n1152, n_2985);
  not g5741 (n_2986, n3396);
  and g5742 (n3397, n1156, n_2986);
  not g5743 (n_2987, n3397);
  and g5744 (n3398, n1160, n_2987);
  not g5745 (n_2988, n3398);
  and g5746 (n3399, n1164, n_2988);
  not g5747 (n_2989, n3399);
  and g5748 (n3400, n1168, n_2989);
  not g5749 (n_2990, n3400);
  and g5750 (n3401, n1172, n_2990);
  not g5751 (n_2991, n3401);
  and g5752 (n3402, n1176, n_2991);
  not g5753 (n_2992, n3402);
  and g5754 (n3403, n1180, n_2992);
  not g5755 (n_2993, n3403);
  and g5756 (n3404, n1184, n_2993);
  not g5757 (n_2994, n3404);
  and g5758 (n3405, n1188, n_2994);
  not g5759 (n_2995, n3405);
  and g5760 (n3406, n1192, n_2995);
  not g5761 (n_2996, n3406);
  and g5762 (n3407, n1196, n_2996);
  not g5763 (n_2997, n3407);
  and g5764 (n3408, n1200, n_2997);
  not g5765 (n_2998, n3408);
  and g5766 (n3409, n1204, n_2998);
  not g5767 (n_2999, n3409);
  and g5768 (n3410, n1208, n_2999);
  not g5769 (n_3000, n3410);
  and g5770 (n3411, n1212, n_3000);
  not g5771 (n_3001, n3411);
  and g5772 (n3412, n1216, n_3001);
  not g5773 (n_3002, n3412);
  and g5774 (n3413, n1220, n_3002);
  not g5775 (n_3003, n3413);
  and g5776 (n3414, n1224, n_3003);
  not g5777 (n_3004, n3414);
  and g5778 (n3415, n1228, n_3004);
  not g5779 (n_3005, n3415);
  and g5780 (n3416, n1232, n_3005);
  not g5781 (n_3006, n3416);
  and g5782 (n3417, n1236, n_3006);
  not g5783 (n_3007, n3417);
  and g5784 (n3418, n1240, n_3007);
  not g5785 (n_3008, n3418);
  and g5786 (n3419, n1244, n_3008);
  not g5787 (n_3009, n3419);
  and g5788 (n3420, n1248, n_3009);
  not g5789 (n_3010, n3420);
  and g5790 (n3421, n1252, n_3010);
  not g5791 (n_3011, n3421);
  and g5792 (n3422, n1256, n_3011);
  not g5793 (n_3012, n3422);
  and g5794 (n3423, n1260, n_3012);
  not g5795 (n_3013, n3423);
  and g5796 (n3424, n1264, n_3013);
  not g5797 (n_3014, n3424);
  and g5798 (n3425, n1268, n_3014);
  not g5799 (n_3015, n3425);
  and g5800 (n3426, n1272, n_3015);
  not g5801 (n_3016, n3426);
  and g5802 (n3427, n1276, n_3016);
  not g5803 (n_3017, n3427);
  and g5804 (n3428, n1280, n_3017);
  not g5805 (n_3018, n3428);
  and g5806 (n3429, n1284, n_3018);
  not g5807 (n_3019, n3429);
  and g5808 (n3430, n1288, n_3019);
  not g5809 (n_3020, n3430);
  and g5810 (n3431, n1292, n_3020);
  not g5811 (n_3021, n3431);
  and g5812 (n3432, n1296, n_3021);
  not g5813 (n_3022, n3432);
  and g5814 (n3433, n1300, n_3022);
  not g5815 (n_3023, n3433);
  and g5816 (n3434, n1304, n_3023);
  not g5817 (n_3024, n3434);
  and g5818 (n3435, n1308, n_3024);
  not g5819 (n_3025, n3435);
  and g5820 (n3436, n1312, n_3025);
  not g5821 (n_3026, n3436);
  and g5822 (n3437, n1316, n_3026);
  not g5823 (n_3027, n3437);
  and g5824 (n3438, n1320, n_3027);
  not g5825 (n_3028, n3438);
  and g5826 (n3439, n1324, n_3028);
  not g5827 (n_3029, n3439);
  and g5828 (n3440, n1328, n_3029);
  not g5829 (n_3030, n3440);
  and g5830 (n3441, n1332, n_3030);
  not g5831 (n_3031, n3441);
  and g5832 (n3442, n1336, n_3031);
  not g5833 (n_3032, n3442);
  and g5834 (n3443, n1340, n_3032);
  not g5835 (n_3033, n3443);
  and g5836 (n3444, n1344, n_3033);
  not g5837 (n_3034, n3444);
  and g5838 (n3445, n1348, n_3034);
  not g5839 (n_3035, n3445);
  and g5840 (n3446, n1352, n_3035);
  not g5841 (n_3036, n3446);
  and g5842 (n3447, n1356, n_3036);
  not g5843 (n_3037, n3447);
  and g5844 (n3448, n1360, n_3037);
  not g5845 (n_3038, n3448);
  and g5846 (n3449, n1364, n_3038);
  not g5847 (n_3039, n3449);
  and g5848 (n3450, n1368, n_3039);
  not g5849 (n_3040, n3450);
  and g5850 (n3451, n1372, n_3040);
  not g5851 (n_3041, n3451);
  and g5852 (n3452, n1376, n_3041);
  not g5853 (n_3042, n3452);
  and g5854 (n3453, n1380, n_3042);
  not g5855 (n_3043, n3453);
  and g5856 (n3454, n1384, n_3043);
  not g5857 (n_3044, n3454);
  and g5858 (n3455, n1388, n_3044);
  not g5859 (n_3045, n3455);
  and g5860 (n3456, n1392, n_3045);
  not g5861 (n_3046, n3456);
  and g5862 (n3457, n1396, n_3046);
  not g5863 (n_3047, n3457);
  and g5864 (n3458, n1663, n_3047);
  not g5865 (n_3048, n3458);
  and g5866 (n3459, n392, n_3048);
  not g5867 (n_3049, n3459);
  and g5868 (n3460, n396, n_3049);
  not g5869 (n_3050, n3460);
  and g5870 (n3461, n400, n_3050);
  not g5871 (n_3051, n3461);
  and g5872 (n3462, n404, n_3051);
  not g5873 (n_3052, n3462);
  and g5874 (n3463, n408, n_3052);
  not g5875 (n_3053, n3463);
  and g5876 (n3464, n412, n_3053);
  not g5877 (n_3054, n3464);
  and g5878 (n3465, n416, n_3054);
  not g5879 (n_3055, n3465);
  and g5880 (n3466, n420, n_3055);
  not g5881 (n_3056, n3466);
  and g5882 (n3467, n424, n_3056);
  not g5883 (n_3057, n3467);
  and g5884 (n3468, n428, n_3057);
  not g5885 (n_3058, n3468);
  and g5886 (n3469, n432, n_3058);
  not g5887 (n_3059, n3469);
  and g5888 (n3470, n436, n_3059);
  not g5889 (n_3060, n3470);
  and g5890 (n3471, n440, n_3060);
  not g5891 (n_3061, n3471);
  and g5892 (n3472, n444, n_3061);
  not g5893 (n_3062, n3472);
  and g5894 (n3473, n448, n_3062);
  and g5895 (n3474, \req[26] , n_122);
  not g5896 (n_3063, n3473);
  and g5897 (\grant[26] , n_3063, n3474);
  not g5898 (n_3064, n794);
  and g5899 (n3476, n459, n_3064);
  not g5900 (n_3065, n3476);
  and g5901 (n3477, n464, n_3065);
  not g5902 (n_3066, n3477);
  and g5903 (n3478, n468, n_3066);
  not g5904 (n_3067, n3478);
  and g5905 (n3479, n472, n_3067);
  not g5906 (n_3068, n3479);
  and g5907 (n3480, n476, n_3068);
  not g5908 (n_3069, n3480);
  and g5909 (n3481, n480, n_3069);
  not g5910 (n_3070, n3481);
  and g5911 (n3482, n484, n_3070);
  not g5912 (n_3071, n3482);
  and g5913 (n3483, n488, n_3071);
  not g5914 (n_3072, n3483);
  and g5915 (n3484, n492, n_3072);
  not g5916 (n_3073, n3484);
  and g5917 (n3485, n496, n_3073);
  not g5918 (n_3074, n3485);
  and g5919 (n3486, n500, n_3074);
  not g5920 (n_3075, n3486);
  and g5921 (n3487, n504, n_3075);
  not g5922 (n_3076, n3487);
  and g5923 (n3488, n508, n_3076);
  not g5924 (n_3077, n3488);
  and g5925 (n3489, n512, n_3077);
  not g5926 (n_3078, n3489);
  and g5927 (n3490, n516, n_3078);
  not g5928 (n_3079, n3490);
  and g5929 (n3491, n520, n_3079);
  not g5930 (n_3080, n3491);
  and g5931 (n3492, n524, n_3080);
  not g5932 (n_3081, n3492);
  and g5933 (n3493, n528, n_3081);
  not g5934 (n_3082, n3493);
  and g5935 (n3494, n532, n_3082);
  not g5936 (n_3083, n3494);
  and g5937 (n3495, n536, n_3083);
  not g5938 (n_3084, n3495);
  and g5939 (n3496, n540, n_3084);
  not g5940 (n_3085, n3496);
  and g5941 (n3497, n544, n_3085);
  not g5942 (n_3086, n3497);
  and g5943 (n3498, n548, n_3086);
  not g5944 (n_3087, n3498);
  and g5945 (n3499, n552, n_3087);
  not g5946 (n_3088, n3499);
  and g5947 (n3500, n556, n_3088);
  not g5948 (n_3089, n3500);
  and g5949 (n3501, n560, n_3089);
  not g5950 (n_3090, n3501);
  and g5951 (n3502, n564, n_3090);
  not g5952 (n_3091, n3502);
  and g5953 (n3503, n568, n_3091);
  not g5954 (n_3092, n3503);
  and g5955 (n3504, n572, n_3092);
  not g5956 (n_3093, n3504);
  and g5957 (n3505, n576, n_3093);
  not g5958 (n_3094, n3505);
  and g5959 (n3506, n580, n_3094);
  not g5960 (n_3095, n3506);
  and g5961 (n3507, n584, n_3095);
  not g5962 (n_3096, n3507);
  and g5963 (n3508, n588, n_3096);
  not g5964 (n_3097, n3508);
  and g5965 (n3509, n592, n_3097);
  not g5966 (n_3098, n3509);
  and g5967 (n3510, n596, n_3098);
  not g5968 (n_3099, n3510);
  and g5969 (n3511, n600, n_3099);
  not g5970 (n_3100, n3511);
  and g5971 (n3512, n604, n_3100);
  not g5972 (n_3101, n3512);
  and g5973 (n3513, n608, n_3101);
  not g5974 (n_3102, n3513);
  and g5975 (n3514, n612, n_3102);
  not g5976 (n_3103, n3514);
  and g5977 (n3515, n616, n_3103);
  not g5978 (n_3104, n3515);
  and g5979 (n3516, n620, n_3104);
  not g5980 (n_3105, n3516);
  and g5981 (n3517, n624, n_3105);
  not g5982 (n_3106, n3517);
  and g5983 (n3518, n628, n_3106);
  not g5984 (n_3107, n3518);
  and g5985 (n3519, n632, n_3107);
  not g5986 (n_3108, n3519);
  and g5987 (n3520, n636, n_3108);
  not g5988 (n_3109, n3520);
  and g5989 (n3521, n640, n_3109);
  not g5990 (n_3110, n3521);
  and g5991 (n3522, n644, n_3110);
  not g5992 (n_3111, n3522);
  and g5993 (n3523, n648, n_3111);
  not g5994 (n_3112, n3523);
  and g5995 (n3524, n652, n_3112);
  not g5996 (n_3113, n3524);
  and g5997 (n3525, n656, n_3113);
  not g5998 (n_3114, n3525);
  and g5999 (n3526, n660, n_3114);
  not g6000 (n_3115, n3526);
  and g6001 (n3527, n664, n_3115);
  not g6002 (n_3116, n3527);
  and g6003 (n3528, n668, n_3116);
  not g6004 (n_3117, n3528);
  and g6005 (n3529, n672, n_3117);
  not g6006 (n_3118, n3529);
  and g6007 (n3530, n676, n_3118);
  not g6008 (n_3119, n3530);
  and g6009 (n3531, n680, n_3119);
  not g6010 (n_3120, n3531);
  and g6011 (n3532, n684, n_3120);
  not g6012 (n_3121, n3532);
  and g6013 (n3533, n688, n_3121);
  not g6014 (n_3122, n3533);
  and g6015 (n3534, n692, n_3122);
  not g6016 (n_3123, n3534);
  and g6017 (n3535, n696, n_3123);
  not g6018 (n_3124, n3535);
  and g6019 (n3536, n700, n_3124);
  not g6020 (n_3125, n3536);
  and g6021 (n3537, n704, n_3125);
  not g6022 (n_3126, n3537);
  and g6023 (n3538, n708, n_3126);
  not g6024 (n_3127, n3538);
  and g6025 (n3539, n712, n_3127);
  not g6026 (n_3128, n3539);
  and g6027 (n3540, n716, n_3128);
  not g6028 (n_3129, n3540);
  and g6029 (n3541, n720, n_3129);
  not g6030 (n_3130, n3541);
  and g6031 (n3542, n1484, n_3130);
  not g6032 (n_3131, n3542);
  and g6033 (n3543, n1486, n_3131);
  not g6034 (n_3132, n3543);
  and g6035 (n3544, n1750, n_3132);
  not g6036 (n_3133, n3544);
  and g6037 (n3545, n731, n_3133);
  not g6038 (n_3134, n3545);
  and g6039 (n3546, n735, n_3134);
  not g6040 (n_3135, n3546);
  and g6041 (n3547, n739, n_3135);
  not g6042 (n_3136, n3547);
  and g6043 (n3548, n743, n_3136);
  not g6044 (n_3137, n3548);
  and g6045 (n3549, n747, n_3137);
  not g6046 (n_3138, n3549);
  and g6047 (n3550, n751, n_3138);
  not g6048 (n_3139, n3550);
  and g6049 (n3551, n755, n_3139);
  not g6050 (n_3140, n3551);
  and g6051 (n3552, n759, n_3140);
  not g6052 (n_3141, n3552);
  and g6053 (n3553, n763, n_3141);
  not g6054 (n_3142, n3553);
  and g6055 (n3554, n767, n_3142);
  not g6056 (n_3143, n3554);
  and g6057 (n3555, n771, n_3143);
  not g6058 (n_3144, n3555);
  and g6059 (n3556, n775, n_3144);
  not g6060 (n_3145, n3556);
  and g6061 (n3557, n779, n_3145);
  not g6062 (n_3146, n3557);
  and g6063 (n3558, n783, n_3146);
  not g6064 (n_3147, n3558);
  and g6065 (n3559, n787, n_3147);
  and g6066 (n3560, \req[27] , n_647);
  not g6067 (n_3148, n3559);
  and g6068 (\grant[27] , n_3148, n3560);
  not g6069 (n_3149, n1131);
  and g6070 (n3562, n798, n_3149);
  not g6071 (n_3150, n3562);
  and g6072 (n3563, n803, n_3150);
  not g6073 (n_3151, n3563);
  and g6074 (n3564, n807, n_3151);
  not g6075 (n_3152, n3564);
  and g6076 (n3565, n811, n_3152);
  not g6077 (n_3153, n3565);
  and g6078 (n3566, n815, n_3153);
  not g6079 (n_3154, n3566);
  and g6080 (n3567, n819, n_3154);
  not g6081 (n_3155, n3567);
  and g6082 (n3568, n823, n_3155);
  not g6083 (n_3156, n3568);
  and g6084 (n3569, n827, n_3156);
  not g6085 (n_3157, n3569);
  and g6086 (n3570, n831, n_3157);
  not g6087 (n_3158, n3570);
  and g6088 (n3571, n835, n_3158);
  not g6089 (n_3159, n3571);
  and g6090 (n3572, n839, n_3159);
  not g6091 (n_3160, n3572);
  and g6092 (n3573, n843, n_3160);
  not g6093 (n_3161, n3573);
  and g6094 (n3574, n847, n_3161);
  not g6095 (n_3162, n3574);
  and g6096 (n3575, n851, n_3162);
  not g6097 (n_3163, n3575);
  and g6098 (n3576, n855, n_3163);
  not g6099 (n_3164, n3576);
  and g6100 (n3577, n859, n_3164);
  not g6101 (n_3165, n3577);
  and g6102 (n3578, n863, n_3165);
  not g6103 (n_3166, n3578);
  and g6104 (n3579, n867, n_3166);
  not g6105 (n_3167, n3579);
  and g6106 (n3580, n871, n_3167);
  not g6107 (n_3168, n3580);
  and g6108 (n3581, n875, n_3168);
  not g6109 (n_3169, n3581);
  and g6110 (n3582, n879, n_3169);
  not g6111 (n_3170, n3582);
  and g6112 (n3583, n883, n_3170);
  not g6113 (n_3171, n3583);
  and g6114 (n3584, n887, n_3171);
  not g6115 (n_3172, n3584);
  and g6116 (n3585, n891, n_3172);
  not g6117 (n_3173, n3585);
  and g6118 (n3586, n895, n_3173);
  not g6119 (n_3174, n3586);
  and g6120 (n3587, n899, n_3174);
  not g6121 (n_3175, n3587);
  and g6122 (n3588, n903, n_3175);
  not g6123 (n_3176, n3588);
  and g6124 (n3589, n907, n_3176);
  not g6125 (n_3177, n3589);
  and g6126 (n3590, n911, n_3177);
  not g6127 (n_3178, n3590);
  and g6128 (n3591, n915, n_3178);
  not g6129 (n_3179, n3591);
  and g6130 (n3592, n919, n_3179);
  not g6131 (n_3180, n3592);
  and g6132 (n3593, n923, n_3180);
  not g6133 (n_3181, n3593);
  and g6134 (n3594, n927, n_3181);
  not g6135 (n_3182, n3594);
  and g6136 (n3595, n931, n_3182);
  not g6137 (n_3183, n3595);
  and g6138 (n3596, n935, n_3183);
  not g6139 (n_3184, n3596);
  and g6140 (n3597, n939, n_3184);
  not g6141 (n_3185, n3597);
  and g6142 (n3598, n943, n_3185);
  not g6143 (n_3186, n3598);
  and g6144 (n3599, n947, n_3186);
  not g6145 (n_3187, n3599);
  and g6146 (n3600, n951, n_3187);
  not g6147 (n_3188, n3600);
  and g6148 (n3601, n955, n_3188);
  not g6149 (n_3189, n3601);
  and g6150 (n3602, n959, n_3189);
  not g6151 (n_3190, n3602);
  and g6152 (n3603, n963, n_3190);
  not g6153 (n_3191, n3603);
  and g6154 (n3604, n967, n_3191);
  not g6155 (n_3192, n3604);
  and g6156 (n3605, n971, n_3192);
  not g6157 (n_3193, n3605);
  and g6158 (n3606, n975, n_3193);
  not g6159 (n_3194, n3606);
  and g6160 (n3607, n979, n_3194);
  not g6161 (n_3195, n3607);
  and g6162 (n3608, n983, n_3195);
  not g6163 (n_3196, n3608);
  and g6164 (n3609, n987, n_3196);
  not g6165 (n_3197, n3609);
  and g6166 (n3610, n991, n_3197);
  not g6167 (n_3198, n3610);
  and g6168 (n3611, n995, n_3198);
  not g6169 (n_3199, n3611);
  and g6170 (n3612, n999, n_3199);
  not g6171 (n_3200, n3612);
  and g6172 (n3613, n1003, n_3200);
  not g6173 (n_3201, n3613);
  and g6174 (n3614, n1007, n_3201);
  not g6175 (n_3202, n3614);
  and g6176 (n3615, n1011, n_3202);
  not g6177 (n_3203, n3615);
  and g6178 (n3616, n1015, n_3203);
  not g6179 (n_3204, n3616);
  and g6180 (n3617, n1019, n_3204);
  not g6181 (n_3205, n3617);
  and g6182 (n3618, n1023, n_3205);
  not g6183 (n_3206, n3618);
  and g6184 (n3619, n1027, n_3206);
  not g6185 (n_3207, n3619);
  and g6186 (n3620, n1031, n_3207);
  not g6187 (n_3208, n3620);
  and g6188 (n3621, n1035, n_3208);
  not g6189 (n_3209, n3621);
  and g6190 (n3622, n1039, n_3209);
  not g6191 (n_3210, n3622);
  and g6192 (n3623, n1043, n_3210);
  not g6193 (n_3211, n3623);
  and g6194 (n3624, n1047, n_3211);
  not g6195 (n_3212, n3624);
  and g6196 (n3625, n1051, n_3212);
  not g6197 (n_3213, n3625);
  and g6198 (n3626, n1055, n_3213);
  not g6199 (n_3214, n3626);
  and g6200 (n3627, n1059, n_3214);
  not g6201 (n_3215, n3627);
  and g6202 (n3628, n1574, n_3215);
  not g6203 (n_3216, n3628);
  and g6204 (n3629, n1576, n_3216);
  not g6205 (n_3217, n3629);
  and g6206 (n3630, n1837, n_3217);
  not g6207 (n_3218, n3630);
  and g6208 (n3631, n1068, n_3218);
  not g6209 (n_3219, n3631);
  and g6210 (n3632, n1072, n_3219);
  not g6211 (n_3220, n3632);
  and g6212 (n3633, n1076, n_3220);
  not g6213 (n_3221, n3633);
  and g6214 (n3634, n1080, n_3221);
  not g6215 (n_3222, n3634);
  and g6216 (n3635, n1084, n_3222);
  not g6217 (n_3223, n3635);
  and g6218 (n3636, n1088, n_3223);
  not g6219 (n_3224, n3636);
  and g6220 (n3637, n1092, n_3224);
  not g6221 (n_3225, n3637);
  and g6222 (n3638, n1096, n_3225);
  not g6223 (n_3226, n3638);
  and g6224 (n3639, n1100, n_3226);
  not g6225 (n_3227, n3639);
  and g6226 (n3640, n1104, n_3227);
  not g6227 (n_3228, n3640);
  and g6228 (n3641, n1108, n_3228);
  not g6229 (n_3229, n3641);
  and g6230 (n3642, n1112, n_3229);
  not g6231 (n_3230, n3642);
  and g6232 (n3643, n1116, n_3230);
  not g6233 (n_3231, n3643);
  and g6234 (n3644, n1120, n_3231);
  not g6235 (n_3232, n3644);
  and g6236 (n3645, n1124, n_3232);
  and g6237 (n3646, \req[28] , n_883);
  not g6238 (n_3233, n3645);
  and g6239 (\grant[28] , n_3233, n3646);
  not g6240 (n_3234, n463);
  and g6241 (n3648, n_3234, n1135);
  not g6242 (n_3235, n3648);
  and g6243 (n3649, n1140, n_3235);
  not g6244 (n_3236, n3649);
  and g6245 (n3650, n1144, n_3236);
  not g6246 (n_3237, n3650);
  and g6247 (n3651, n1148, n_3237);
  not g6248 (n_3238, n3651);
  and g6249 (n3652, n1152, n_3238);
  not g6250 (n_3239, n3652);
  and g6251 (n3653, n1156, n_3239);
  not g6252 (n_3240, n3653);
  and g6253 (n3654, n1160, n_3240);
  not g6254 (n_3241, n3654);
  and g6255 (n3655, n1164, n_3241);
  not g6256 (n_3242, n3655);
  and g6257 (n3656, n1168, n_3242);
  not g6258 (n_3243, n3656);
  and g6259 (n3657, n1172, n_3243);
  not g6260 (n_3244, n3657);
  and g6261 (n3658, n1176, n_3244);
  not g6262 (n_3245, n3658);
  and g6263 (n3659, n1180, n_3245);
  not g6264 (n_3246, n3659);
  and g6265 (n3660, n1184, n_3246);
  not g6266 (n_3247, n3660);
  and g6267 (n3661, n1188, n_3247);
  not g6268 (n_3248, n3661);
  and g6269 (n3662, n1192, n_3248);
  not g6270 (n_3249, n3662);
  and g6271 (n3663, n1196, n_3249);
  not g6272 (n_3250, n3663);
  and g6273 (n3664, n1200, n_3250);
  not g6274 (n_3251, n3664);
  and g6275 (n3665, n1204, n_3251);
  not g6276 (n_3252, n3665);
  and g6277 (n3666, n1208, n_3252);
  not g6278 (n_3253, n3666);
  and g6279 (n3667, n1212, n_3253);
  not g6280 (n_3254, n3667);
  and g6281 (n3668, n1216, n_3254);
  not g6282 (n_3255, n3668);
  and g6283 (n3669, n1220, n_3255);
  not g6284 (n_3256, n3669);
  and g6285 (n3670, n1224, n_3256);
  not g6286 (n_3257, n3670);
  and g6287 (n3671, n1228, n_3257);
  not g6288 (n_3258, n3671);
  and g6289 (n3672, n1232, n_3258);
  not g6290 (n_3259, n3672);
  and g6291 (n3673, n1236, n_3259);
  not g6292 (n_3260, n3673);
  and g6293 (n3674, n1240, n_3260);
  not g6294 (n_3261, n3674);
  and g6295 (n3675, n1244, n_3261);
  not g6296 (n_3262, n3675);
  and g6297 (n3676, n1248, n_3262);
  not g6298 (n_3263, n3676);
  and g6299 (n3677, n1252, n_3263);
  not g6300 (n_3264, n3677);
  and g6301 (n3678, n1256, n_3264);
  not g6302 (n_3265, n3678);
  and g6303 (n3679, n1260, n_3265);
  not g6304 (n_3266, n3679);
  and g6305 (n3680, n1264, n_3266);
  not g6306 (n_3267, n3680);
  and g6307 (n3681, n1268, n_3267);
  not g6308 (n_3268, n3681);
  and g6309 (n3682, n1272, n_3268);
  not g6310 (n_3269, n3682);
  and g6311 (n3683, n1276, n_3269);
  not g6312 (n_3270, n3683);
  and g6313 (n3684, n1280, n_3270);
  not g6314 (n_3271, n3684);
  and g6315 (n3685, n1284, n_3271);
  not g6316 (n_3272, n3685);
  and g6317 (n3686, n1288, n_3272);
  not g6318 (n_3273, n3686);
  and g6319 (n3687, n1292, n_3273);
  not g6320 (n_3274, n3687);
  and g6321 (n3688, n1296, n_3274);
  not g6322 (n_3275, n3688);
  and g6323 (n3689, n1300, n_3275);
  not g6324 (n_3276, n3689);
  and g6325 (n3690, n1304, n_3276);
  not g6326 (n_3277, n3690);
  and g6327 (n3691, n1308, n_3277);
  not g6328 (n_3278, n3691);
  and g6329 (n3692, n1312, n_3278);
  not g6330 (n_3279, n3692);
  and g6331 (n3693, n1316, n_3279);
  not g6332 (n_3280, n3693);
  and g6333 (n3694, n1320, n_3280);
  not g6334 (n_3281, n3694);
  and g6335 (n3695, n1324, n_3281);
  not g6336 (n_3282, n3695);
  and g6337 (n3696, n1328, n_3282);
  not g6338 (n_3283, n3696);
  and g6339 (n3697, n1332, n_3283);
  not g6340 (n_3284, n3697);
  and g6341 (n3698, n1336, n_3284);
  not g6342 (n_3285, n3698);
  and g6343 (n3699, n1340, n_3285);
  not g6344 (n_3286, n3699);
  and g6345 (n3700, n1344, n_3286);
  not g6346 (n_3287, n3700);
  and g6347 (n3701, n1348, n_3287);
  not g6348 (n_3288, n3701);
  and g6349 (n3702, n1352, n_3288);
  not g6350 (n_3289, n3702);
  and g6351 (n3703, n1356, n_3289);
  not g6352 (n_3290, n3703);
  and g6353 (n3704, n1360, n_3290);
  not g6354 (n_3291, n3704);
  and g6355 (n3705, n1364, n_3291);
  not g6356 (n_3292, n3705);
  and g6357 (n3706, n1368, n_3292);
  not g6358 (n_3293, n3706);
  and g6359 (n3707, n1372, n_3293);
  not g6360 (n_3294, n3707);
  and g6361 (n3708, n1376, n_3294);
  not g6362 (n_3295, n3708);
  and g6363 (n3709, n1380, n_3295);
  not g6364 (n_3296, n3709);
  and g6365 (n3710, n1384, n_3296);
  not g6366 (n_3297, n3710);
  and g6367 (n3711, n1388, n_3297);
  not g6368 (n_3298, n3711);
  and g6369 (n3712, n1392, n_3298);
  not g6370 (n_3299, n3712);
  and g6371 (n3713, n1396, n_3299);
  not g6372 (n_3300, n3713);
  and g6373 (n3714, n1663, n_3300);
  not g6374 (n_3301, n3714);
  and g6375 (n3715, n392, n_3301);
  not g6376 (n_3302, n3715);
  and g6377 (n3716, n396, n_3302);
  not g6378 (n_3303, n3716);
  and g6379 (n3717, n400, n_3303);
  not g6380 (n_3304, n3717);
  and g6381 (n3718, n404, n_3304);
  not g6382 (n_3305, n3718);
  and g6383 (n3719, n408, n_3305);
  not g6384 (n_3306, n3719);
  and g6385 (n3720, n412, n_3306);
  not g6386 (n_3307, n3720);
  and g6387 (n3721, n416, n_3307);
  not g6388 (n_3308, n3721);
  and g6389 (n3722, n420, n_3308);
  not g6390 (n_3309, n3722);
  and g6391 (n3723, n424, n_3309);
  not g6392 (n_3310, n3723);
  and g6393 (n3724, n428, n_3310);
  not g6394 (n_3311, n3724);
  and g6395 (n3725, n432, n_3311);
  not g6396 (n_3312, n3725);
  and g6397 (n3726, n436, n_3312);
  not g6398 (n_3313, n3726);
  and g6399 (n3727, n440, n_3313);
  not g6400 (n_3314, n3727);
  and g6401 (n3728, n444, n_3314);
  not g6402 (n_3315, n3728);
  and g6403 (n3729, n448, n_3315);
  not g6404 (n_3316, n3729);
  and g6405 (n3730, n452, n_3316);
  not g6406 (n_3317, n3730);
  and g6407 (n3731, n456, n_3317);
  and g6408 (n3732, \req[29] , n_136);
  not g6409 (n_3318, n3731);
  and g6410 (\grant[29] , n_3318, n3732);
  not g6411 (n_3319, n802);
  and g6412 (n3734, n467, n_3319);
  not g6413 (n_3320, n3734);
  and g6414 (n3735, n472, n_3320);
  not g6415 (n_3321, n3735);
  and g6416 (n3736, n476, n_3321);
  not g6417 (n_3322, n3736);
  and g6418 (n3737, n480, n_3322);
  not g6419 (n_3323, n3737);
  and g6420 (n3738, n484, n_3323);
  not g6421 (n_3324, n3738);
  and g6422 (n3739, n488, n_3324);
  not g6423 (n_3325, n3739);
  and g6424 (n3740, n492, n_3325);
  not g6425 (n_3326, n3740);
  and g6426 (n3741, n496, n_3326);
  not g6427 (n_3327, n3741);
  and g6428 (n3742, n500, n_3327);
  not g6429 (n_3328, n3742);
  and g6430 (n3743, n504, n_3328);
  not g6431 (n_3329, n3743);
  and g6432 (n3744, n508, n_3329);
  not g6433 (n_3330, n3744);
  and g6434 (n3745, n512, n_3330);
  not g6435 (n_3331, n3745);
  and g6436 (n3746, n516, n_3331);
  not g6437 (n_3332, n3746);
  and g6438 (n3747, n520, n_3332);
  not g6439 (n_3333, n3747);
  and g6440 (n3748, n524, n_3333);
  not g6441 (n_3334, n3748);
  and g6442 (n3749, n528, n_3334);
  not g6443 (n_3335, n3749);
  and g6444 (n3750, n532, n_3335);
  not g6445 (n_3336, n3750);
  and g6446 (n3751, n536, n_3336);
  not g6447 (n_3337, n3751);
  and g6448 (n3752, n540, n_3337);
  not g6449 (n_3338, n3752);
  and g6450 (n3753, n544, n_3338);
  not g6451 (n_3339, n3753);
  and g6452 (n3754, n548, n_3339);
  not g6453 (n_3340, n3754);
  and g6454 (n3755, n552, n_3340);
  not g6455 (n_3341, n3755);
  and g6456 (n3756, n556, n_3341);
  not g6457 (n_3342, n3756);
  and g6458 (n3757, n560, n_3342);
  not g6459 (n_3343, n3757);
  and g6460 (n3758, n564, n_3343);
  not g6461 (n_3344, n3758);
  and g6462 (n3759, n568, n_3344);
  not g6463 (n_3345, n3759);
  and g6464 (n3760, n572, n_3345);
  not g6465 (n_3346, n3760);
  and g6466 (n3761, n576, n_3346);
  not g6467 (n_3347, n3761);
  and g6468 (n3762, n580, n_3347);
  not g6469 (n_3348, n3762);
  and g6470 (n3763, n584, n_3348);
  not g6471 (n_3349, n3763);
  and g6472 (n3764, n588, n_3349);
  not g6473 (n_3350, n3764);
  and g6474 (n3765, n592, n_3350);
  not g6475 (n_3351, n3765);
  and g6476 (n3766, n596, n_3351);
  not g6477 (n_3352, n3766);
  and g6478 (n3767, n600, n_3352);
  not g6479 (n_3353, n3767);
  and g6480 (n3768, n604, n_3353);
  not g6481 (n_3354, n3768);
  and g6482 (n3769, n608, n_3354);
  not g6483 (n_3355, n3769);
  and g6484 (n3770, n612, n_3355);
  not g6485 (n_3356, n3770);
  and g6486 (n3771, n616, n_3356);
  not g6487 (n_3357, n3771);
  and g6488 (n3772, n620, n_3357);
  not g6489 (n_3358, n3772);
  and g6490 (n3773, n624, n_3358);
  not g6491 (n_3359, n3773);
  and g6492 (n3774, n628, n_3359);
  not g6493 (n_3360, n3774);
  and g6494 (n3775, n632, n_3360);
  not g6495 (n_3361, n3775);
  and g6496 (n3776, n636, n_3361);
  not g6497 (n_3362, n3776);
  and g6498 (n3777, n640, n_3362);
  not g6499 (n_3363, n3777);
  and g6500 (n3778, n644, n_3363);
  not g6501 (n_3364, n3778);
  and g6502 (n3779, n648, n_3364);
  not g6503 (n_3365, n3779);
  and g6504 (n3780, n652, n_3365);
  not g6505 (n_3366, n3780);
  and g6506 (n3781, n656, n_3366);
  not g6507 (n_3367, n3781);
  and g6508 (n3782, n660, n_3367);
  not g6509 (n_3368, n3782);
  and g6510 (n3783, n664, n_3368);
  not g6511 (n_3369, n3783);
  and g6512 (n3784, n668, n_3369);
  not g6513 (n_3370, n3784);
  and g6514 (n3785, n672, n_3370);
  not g6515 (n_3371, n3785);
  and g6516 (n3786, n676, n_3371);
  not g6517 (n_3372, n3786);
  and g6518 (n3787, n680, n_3372);
  not g6519 (n_3373, n3787);
  and g6520 (n3788, n684, n_3373);
  not g6521 (n_3374, n3788);
  and g6522 (n3789, n688, n_3374);
  not g6523 (n_3375, n3789);
  and g6524 (n3790, n692, n_3375);
  not g6525 (n_3376, n3790);
  and g6526 (n3791, n696, n_3376);
  not g6527 (n_3377, n3791);
  and g6528 (n3792, n700, n_3377);
  not g6529 (n_3378, n3792);
  and g6530 (n3793, n704, n_3378);
  not g6531 (n_3379, n3793);
  and g6532 (n3794, n708, n_3379);
  not g6533 (n_3380, n3794);
  and g6534 (n3795, n712, n_3380);
  not g6535 (n_3381, n3795);
  and g6536 (n3796, n716, n_3381);
  not g6537 (n_3382, n3796);
  and g6538 (n3797, n720, n_3382);
  not g6539 (n_3383, n3797);
  and g6540 (n3798, n1484, n_3383);
  not g6541 (n_3384, n3798);
  and g6542 (n3799, n1486, n_3384);
  not g6543 (n_3385, n3799);
  and g6544 (n3800, n1750, n_3385);
  not g6545 (n_3386, n3800);
  and g6546 (n3801, n731, n_3386);
  not g6547 (n_3387, n3801);
  and g6548 (n3802, n735, n_3387);
  not g6549 (n_3388, n3802);
  and g6550 (n3803, n739, n_3388);
  not g6551 (n_3389, n3803);
  and g6552 (n3804, n743, n_3389);
  not g6553 (n_3390, n3804);
  and g6554 (n3805, n747, n_3390);
  not g6555 (n_3391, n3805);
  and g6556 (n3806, n751, n_3391);
  not g6557 (n_3392, n3806);
  and g6558 (n3807, n755, n_3392);
  not g6559 (n_3393, n3807);
  and g6560 (n3808, n759, n_3393);
  not g6561 (n_3394, n3808);
  and g6562 (n3809, n763, n_3394);
  not g6563 (n_3395, n3809);
  and g6564 (n3810, n767, n_3395);
  not g6565 (n_3396, n3810);
  and g6566 (n3811, n771, n_3396);
  not g6567 (n_3397, n3811);
  and g6568 (n3812, n775, n_3397);
  not g6569 (n_3398, n3812);
  and g6570 (n3813, n779, n_3398);
  not g6571 (n_3399, n3813);
  and g6572 (n3814, n783, n_3399);
  not g6573 (n_3400, n3814);
  and g6574 (n3815, n787, n_3400);
  not g6575 (n_3401, n3815);
  and g6576 (n3816, n791, n_3401);
  not g6577 (n_3402, n3816);
  and g6578 (n3817, n795, n_3402);
  and g6579 (n3818, \req[30] , n_653);
  not g6580 (n_3403, n3817);
  and g6581 (\grant[30] , n_3403, n3818);
  not g6582 (n_3404, n1139);
  and g6583 (n3820, n806, n_3404);
  not g6584 (n_3405, n3820);
  and g6585 (n3821, n811, n_3405);
  not g6586 (n_3406, n3821);
  and g6587 (n3822, n815, n_3406);
  not g6588 (n_3407, n3822);
  and g6589 (n3823, n819, n_3407);
  not g6590 (n_3408, n3823);
  and g6591 (n3824, n823, n_3408);
  not g6592 (n_3409, n3824);
  and g6593 (n3825, n827, n_3409);
  not g6594 (n_3410, n3825);
  and g6595 (n3826, n831, n_3410);
  not g6596 (n_3411, n3826);
  and g6597 (n3827, n835, n_3411);
  not g6598 (n_3412, n3827);
  and g6599 (n3828, n839, n_3412);
  not g6600 (n_3413, n3828);
  and g6601 (n3829, n843, n_3413);
  not g6602 (n_3414, n3829);
  and g6603 (n3830, n847, n_3414);
  not g6604 (n_3415, n3830);
  and g6605 (n3831, n851, n_3415);
  not g6606 (n_3416, n3831);
  and g6607 (n3832, n855, n_3416);
  not g6608 (n_3417, n3832);
  and g6609 (n3833, n859, n_3417);
  not g6610 (n_3418, n3833);
  and g6611 (n3834, n863, n_3418);
  not g6612 (n_3419, n3834);
  and g6613 (n3835, n867, n_3419);
  not g6614 (n_3420, n3835);
  and g6615 (n3836, n871, n_3420);
  not g6616 (n_3421, n3836);
  and g6617 (n3837, n875, n_3421);
  not g6618 (n_3422, n3837);
  and g6619 (n3838, n879, n_3422);
  not g6620 (n_3423, n3838);
  and g6621 (n3839, n883, n_3423);
  not g6622 (n_3424, n3839);
  and g6623 (n3840, n887, n_3424);
  not g6624 (n_3425, n3840);
  and g6625 (n3841, n891, n_3425);
  not g6626 (n_3426, n3841);
  and g6627 (n3842, n895, n_3426);
  not g6628 (n_3427, n3842);
  and g6629 (n3843, n899, n_3427);
  not g6630 (n_3428, n3843);
  and g6631 (n3844, n903, n_3428);
  not g6632 (n_3429, n3844);
  and g6633 (n3845, n907, n_3429);
  not g6634 (n_3430, n3845);
  and g6635 (n3846, n911, n_3430);
  not g6636 (n_3431, n3846);
  and g6637 (n3847, n915, n_3431);
  not g6638 (n_3432, n3847);
  and g6639 (n3848, n919, n_3432);
  not g6640 (n_3433, n3848);
  and g6641 (n3849, n923, n_3433);
  not g6642 (n_3434, n3849);
  and g6643 (n3850, n927, n_3434);
  not g6644 (n_3435, n3850);
  and g6645 (n3851, n931, n_3435);
  not g6646 (n_3436, n3851);
  and g6647 (n3852, n935, n_3436);
  not g6648 (n_3437, n3852);
  and g6649 (n3853, n939, n_3437);
  not g6650 (n_3438, n3853);
  and g6651 (n3854, n943, n_3438);
  not g6652 (n_3439, n3854);
  and g6653 (n3855, n947, n_3439);
  not g6654 (n_3440, n3855);
  and g6655 (n3856, n951, n_3440);
  not g6656 (n_3441, n3856);
  and g6657 (n3857, n955, n_3441);
  not g6658 (n_3442, n3857);
  and g6659 (n3858, n959, n_3442);
  not g6660 (n_3443, n3858);
  and g6661 (n3859, n963, n_3443);
  not g6662 (n_3444, n3859);
  and g6663 (n3860, n967, n_3444);
  not g6664 (n_3445, n3860);
  and g6665 (n3861, n971, n_3445);
  not g6666 (n_3446, n3861);
  and g6667 (n3862, n975, n_3446);
  not g6668 (n_3447, n3862);
  and g6669 (n3863, n979, n_3447);
  not g6670 (n_3448, n3863);
  and g6671 (n3864, n983, n_3448);
  not g6672 (n_3449, n3864);
  and g6673 (n3865, n987, n_3449);
  not g6674 (n_3450, n3865);
  and g6675 (n3866, n991, n_3450);
  not g6676 (n_3451, n3866);
  and g6677 (n3867, n995, n_3451);
  not g6678 (n_3452, n3867);
  and g6679 (n3868, n999, n_3452);
  not g6680 (n_3453, n3868);
  and g6681 (n3869, n1003, n_3453);
  not g6682 (n_3454, n3869);
  and g6683 (n3870, n1007, n_3454);
  not g6684 (n_3455, n3870);
  and g6685 (n3871, n1011, n_3455);
  not g6686 (n_3456, n3871);
  and g6687 (n3872, n1015, n_3456);
  not g6688 (n_3457, n3872);
  and g6689 (n3873, n1019, n_3457);
  not g6690 (n_3458, n3873);
  and g6691 (n3874, n1023, n_3458);
  not g6692 (n_3459, n3874);
  and g6693 (n3875, n1027, n_3459);
  not g6694 (n_3460, n3875);
  and g6695 (n3876, n1031, n_3460);
  not g6696 (n_3461, n3876);
  and g6697 (n3877, n1035, n_3461);
  not g6698 (n_3462, n3877);
  and g6699 (n3878, n1039, n_3462);
  not g6700 (n_3463, n3878);
  and g6701 (n3879, n1043, n_3463);
  not g6702 (n_3464, n3879);
  and g6703 (n3880, n1047, n_3464);
  not g6704 (n_3465, n3880);
  and g6705 (n3881, n1051, n_3465);
  not g6706 (n_3466, n3881);
  and g6707 (n3882, n1055, n_3466);
  not g6708 (n_3467, n3882);
  and g6709 (n3883, n1059, n_3467);
  not g6710 (n_3468, n3883);
  and g6711 (n3884, n1574, n_3468);
  not g6712 (n_3469, n3884);
  and g6713 (n3885, n1576, n_3469);
  not g6714 (n_3470, n3885);
  and g6715 (n3886, n1837, n_3470);
  not g6716 (n_3471, n3886);
  and g6717 (n3887, n1068, n_3471);
  not g6718 (n_3472, n3887);
  and g6719 (n3888, n1072, n_3472);
  not g6720 (n_3473, n3888);
  and g6721 (n3889, n1076, n_3473);
  not g6722 (n_3474, n3889);
  and g6723 (n3890, n1080, n_3474);
  not g6724 (n_3475, n3890);
  and g6725 (n3891, n1084, n_3475);
  not g6726 (n_3476, n3891);
  and g6727 (n3892, n1088, n_3476);
  not g6728 (n_3477, n3892);
  and g6729 (n3893, n1092, n_3477);
  not g6730 (n_3478, n3893);
  and g6731 (n3894, n1096, n_3478);
  not g6732 (n_3479, n3894);
  and g6733 (n3895, n1100, n_3479);
  not g6734 (n_3480, n3895);
  and g6735 (n3896, n1104, n_3480);
  not g6736 (n_3481, n3896);
  and g6737 (n3897, n1108, n_3481);
  not g6738 (n_3482, n3897);
  and g6739 (n3898, n1112, n_3482);
  not g6740 (n_3483, n3898);
  and g6741 (n3899, n1116, n_3483);
  not g6742 (n_3484, n3899);
  and g6743 (n3900, n1120, n_3484);
  not g6744 (n_3485, n3900);
  and g6745 (n3901, n1124, n_3485);
  not g6746 (n_3486, n3901);
  and g6747 (n3902, n1128, n_3486);
  not g6748 (n_3487, n3902);
  and g6749 (n3903, n1132, n_3487);
  and g6750 (n3904, \req[31] , n_887);
  not g6751 (n_3488, n3903);
  and g6752 (\grant[31] , n_3488, n3904);
  not g6753 (n_3489, n471);
  and g6754 (n3906, n_3489, n1143);
  not g6755 (n_3490, n3906);
  and g6756 (n3907, n1148, n_3490);
  not g6757 (n_3491, n3907);
  and g6758 (n3908, n1152, n_3491);
  not g6759 (n_3492, n3908);
  and g6760 (n3909, n1156, n_3492);
  not g6761 (n_3493, n3909);
  and g6762 (n3910, n1160, n_3493);
  not g6763 (n_3494, n3910);
  and g6764 (n3911, n1164, n_3494);
  not g6765 (n_3495, n3911);
  and g6766 (n3912, n1168, n_3495);
  not g6767 (n_3496, n3912);
  and g6768 (n3913, n1172, n_3496);
  not g6769 (n_3497, n3913);
  and g6770 (n3914, n1176, n_3497);
  not g6771 (n_3498, n3914);
  and g6772 (n3915, n1180, n_3498);
  not g6773 (n_3499, n3915);
  and g6774 (n3916, n1184, n_3499);
  not g6775 (n_3500, n3916);
  and g6776 (n3917, n1188, n_3500);
  not g6777 (n_3501, n3917);
  and g6778 (n3918, n1192, n_3501);
  not g6779 (n_3502, n3918);
  and g6780 (n3919, n1196, n_3502);
  not g6781 (n_3503, n3919);
  and g6782 (n3920, n1200, n_3503);
  not g6783 (n_3504, n3920);
  and g6784 (n3921, n1204, n_3504);
  not g6785 (n_3505, n3921);
  and g6786 (n3922, n1208, n_3505);
  not g6787 (n_3506, n3922);
  and g6788 (n3923, n1212, n_3506);
  not g6789 (n_3507, n3923);
  and g6790 (n3924, n1216, n_3507);
  not g6791 (n_3508, n3924);
  and g6792 (n3925, n1220, n_3508);
  not g6793 (n_3509, n3925);
  and g6794 (n3926, n1224, n_3509);
  not g6795 (n_3510, n3926);
  and g6796 (n3927, n1228, n_3510);
  not g6797 (n_3511, n3927);
  and g6798 (n3928, n1232, n_3511);
  not g6799 (n_3512, n3928);
  and g6800 (n3929, n1236, n_3512);
  not g6801 (n_3513, n3929);
  and g6802 (n3930, n1240, n_3513);
  not g6803 (n_3514, n3930);
  and g6804 (n3931, n1244, n_3514);
  not g6805 (n_3515, n3931);
  and g6806 (n3932, n1248, n_3515);
  not g6807 (n_3516, n3932);
  and g6808 (n3933, n1252, n_3516);
  not g6809 (n_3517, n3933);
  and g6810 (n3934, n1256, n_3517);
  not g6811 (n_3518, n3934);
  and g6812 (n3935, n1260, n_3518);
  not g6813 (n_3519, n3935);
  and g6814 (n3936, n1264, n_3519);
  not g6815 (n_3520, n3936);
  and g6816 (n3937, n1268, n_3520);
  not g6817 (n_3521, n3937);
  and g6818 (n3938, n1272, n_3521);
  not g6819 (n_3522, n3938);
  and g6820 (n3939, n1276, n_3522);
  not g6821 (n_3523, n3939);
  and g6822 (n3940, n1280, n_3523);
  not g6823 (n_3524, n3940);
  and g6824 (n3941, n1284, n_3524);
  not g6825 (n_3525, n3941);
  and g6826 (n3942, n1288, n_3525);
  not g6827 (n_3526, n3942);
  and g6828 (n3943, n1292, n_3526);
  not g6829 (n_3527, n3943);
  and g6830 (n3944, n1296, n_3527);
  not g6831 (n_3528, n3944);
  and g6832 (n3945, n1300, n_3528);
  not g6833 (n_3529, n3945);
  and g6834 (n3946, n1304, n_3529);
  not g6835 (n_3530, n3946);
  and g6836 (n3947, n1308, n_3530);
  not g6837 (n_3531, n3947);
  and g6838 (n3948, n1312, n_3531);
  not g6839 (n_3532, n3948);
  and g6840 (n3949, n1316, n_3532);
  not g6841 (n_3533, n3949);
  and g6842 (n3950, n1320, n_3533);
  not g6843 (n_3534, n3950);
  and g6844 (n3951, n1324, n_3534);
  not g6845 (n_3535, n3951);
  and g6846 (n3952, n1328, n_3535);
  not g6847 (n_3536, n3952);
  and g6848 (n3953, n1332, n_3536);
  not g6849 (n_3537, n3953);
  and g6850 (n3954, n1336, n_3537);
  not g6851 (n_3538, n3954);
  and g6852 (n3955, n1340, n_3538);
  not g6853 (n_3539, n3955);
  and g6854 (n3956, n1344, n_3539);
  not g6855 (n_3540, n3956);
  and g6856 (n3957, n1348, n_3540);
  not g6857 (n_3541, n3957);
  and g6858 (n3958, n1352, n_3541);
  not g6859 (n_3542, n3958);
  and g6860 (n3959, n1356, n_3542);
  not g6861 (n_3543, n3959);
  and g6862 (n3960, n1360, n_3543);
  not g6863 (n_3544, n3960);
  and g6864 (n3961, n1364, n_3544);
  not g6865 (n_3545, n3961);
  and g6866 (n3962, n1368, n_3545);
  not g6867 (n_3546, n3962);
  and g6868 (n3963, n1372, n_3546);
  not g6869 (n_3547, n3963);
  and g6870 (n3964, n1376, n_3547);
  not g6871 (n_3548, n3964);
  and g6872 (n3965, n1380, n_3548);
  not g6873 (n_3549, n3965);
  and g6874 (n3966, n1384, n_3549);
  not g6875 (n_3550, n3966);
  and g6876 (n3967, n1388, n_3550);
  not g6877 (n_3551, n3967);
  and g6878 (n3968, n1392, n_3551);
  not g6879 (n_3552, n3968);
  and g6880 (n3969, n1396, n_3552);
  not g6881 (n_3553, n3969);
  and g6882 (n3970, n1663, n_3553);
  not g6883 (n_3554, n3970);
  and g6884 (n3971, n392, n_3554);
  not g6885 (n_3555, n3971);
  and g6886 (n3972, n396, n_3555);
  not g6887 (n_3556, n3972);
  and g6888 (n3973, n400, n_3556);
  not g6889 (n_3557, n3973);
  and g6890 (n3974, n404, n_3557);
  not g6891 (n_3558, n3974);
  and g6892 (n3975, n408, n_3558);
  not g6893 (n_3559, n3975);
  and g6894 (n3976, n412, n_3559);
  not g6895 (n_3560, n3976);
  and g6896 (n3977, n416, n_3560);
  not g6897 (n_3561, n3977);
  and g6898 (n3978, n420, n_3561);
  not g6899 (n_3562, n3978);
  and g6900 (n3979, n424, n_3562);
  not g6901 (n_3563, n3979);
  and g6902 (n3980, n428, n_3563);
  not g6903 (n_3564, n3980);
  and g6904 (n3981, n432, n_3564);
  not g6905 (n_3565, n3981);
  and g6906 (n3982, n436, n_3565);
  not g6907 (n_3566, n3982);
  and g6908 (n3983, n440, n_3566);
  not g6909 (n_3567, n3983);
  and g6910 (n3984, n444, n_3567);
  not g6911 (n_3568, n3984);
  and g6912 (n3985, n448, n_3568);
  not g6913 (n_3569, n3985);
  and g6914 (n3986, n452, n_3569);
  not g6915 (n_3570, n3986);
  and g6916 (n3987, n456, n_3570);
  not g6917 (n_3571, n3987);
  and g6918 (n3988, n460, n_3571);
  not g6919 (n_3572, n3988);
  and g6920 (n3989, n464, n_3572);
  and g6921 (n3990, \req[32] , n_150);
  not g6922 (n_3573, n3989);
  and g6923 (\grant[32] , n_3573, n3990);
  not g6924 (n_3574, n810);
  and g6925 (n3992, n475, n_3574);
  not g6926 (n_3575, n3992);
  and g6927 (n3993, n480, n_3575);
  not g6928 (n_3576, n3993);
  and g6929 (n3994, n484, n_3576);
  not g6930 (n_3577, n3994);
  and g6931 (n3995, n488, n_3577);
  not g6932 (n_3578, n3995);
  and g6933 (n3996, n492, n_3578);
  not g6934 (n_3579, n3996);
  and g6935 (n3997, n496, n_3579);
  not g6936 (n_3580, n3997);
  and g6937 (n3998, n500, n_3580);
  not g6938 (n_3581, n3998);
  and g6939 (n3999, n504, n_3581);
  not g6940 (n_3582, n3999);
  and g6941 (n4000, n508, n_3582);
  not g6942 (n_3583, n4000);
  and g6943 (n4001, n512, n_3583);
  not g6944 (n_3584, n4001);
  and g6945 (n4002, n516, n_3584);
  not g6946 (n_3585, n4002);
  and g6947 (n4003, n520, n_3585);
  not g6948 (n_3586, n4003);
  and g6949 (n4004, n524, n_3586);
  not g6950 (n_3587, n4004);
  and g6951 (n4005, n528, n_3587);
  not g6952 (n_3588, n4005);
  and g6953 (n4006, n532, n_3588);
  not g6954 (n_3589, n4006);
  and g6955 (n4007, n536, n_3589);
  not g6956 (n_3590, n4007);
  and g6957 (n4008, n540, n_3590);
  not g6958 (n_3591, n4008);
  and g6959 (n4009, n544, n_3591);
  not g6960 (n_3592, n4009);
  and g6961 (n4010, n548, n_3592);
  not g6962 (n_3593, n4010);
  and g6963 (n4011, n552, n_3593);
  not g6964 (n_3594, n4011);
  and g6965 (n4012, n556, n_3594);
  not g6966 (n_3595, n4012);
  and g6967 (n4013, n560, n_3595);
  not g6968 (n_3596, n4013);
  and g6969 (n4014, n564, n_3596);
  not g6970 (n_3597, n4014);
  and g6971 (n4015, n568, n_3597);
  not g6972 (n_3598, n4015);
  and g6973 (n4016, n572, n_3598);
  not g6974 (n_3599, n4016);
  and g6975 (n4017, n576, n_3599);
  not g6976 (n_3600, n4017);
  and g6977 (n4018, n580, n_3600);
  not g6978 (n_3601, n4018);
  and g6979 (n4019, n584, n_3601);
  not g6980 (n_3602, n4019);
  and g6981 (n4020, n588, n_3602);
  not g6982 (n_3603, n4020);
  and g6983 (n4021, n592, n_3603);
  not g6984 (n_3604, n4021);
  and g6985 (n4022, n596, n_3604);
  not g6986 (n_3605, n4022);
  and g6987 (n4023, n600, n_3605);
  not g6988 (n_3606, n4023);
  and g6989 (n4024, n604, n_3606);
  not g6990 (n_3607, n4024);
  and g6991 (n4025, n608, n_3607);
  not g6992 (n_3608, n4025);
  and g6993 (n4026, n612, n_3608);
  not g6994 (n_3609, n4026);
  and g6995 (n4027, n616, n_3609);
  not g6996 (n_3610, n4027);
  and g6997 (n4028, n620, n_3610);
  not g6998 (n_3611, n4028);
  and g6999 (n4029, n624, n_3611);
  not g7000 (n_3612, n4029);
  and g7001 (n4030, n628, n_3612);
  not g7002 (n_3613, n4030);
  and g7003 (n4031, n632, n_3613);
  not g7004 (n_3614, n4031);
  and g7005 (n4032, n636, n_3614);
  not g7006 (n_3615, n4032);
  and g7007 (n4033, n640, n_3615);
  not g7008 (n_3616, n4033);
  and g7009 (n4034, n644, n_3616);
  not g7010 (n_3617, n4034);
  and g7011 (n4035, n648, n_3617);
  not g7012 (n_3618, n4035);
  and g7013 (n4036, n652, n_3618);
  not g7014 (n_3619, n4036);
  and g7015 (n4037, n656, n_3619);
  not g7016 (n_3620, n4037);
  and g7017 (n4038, n660, n_3620);
  not g7018 (n_3621, n4038);
  and g7019 (n4039, n664, n_3621);
  not g7020 (n_3622, n4039);
  and g7021 (n4040, n668, n_3622);
  not g7022 (n_3623, n4040);
  and g7023 (n4041, n672, n_3623);
  not g7024 (n_3624, n4041);
  and g7025 (n4042, n676, n_3624);
  not g7026 (n_3625, n4042);
  and g7027 (n4043, n680, n_3625);
  not g7028 (n_3626, n4043);
  and g7029 (n4044, n684, n_3626);
  not g7030 (n_3627, n4044);
  and g7031 (n4045, n688, n_3627);
  not g7032 (n_3628, n4045);
  and g7033 (n4046, n692, n_3628);
  not g7034 (n_3629, n4046);
  and g7035 (n4047, n696, n_3629);
  not g7036 (n_3630, n4047);
  and g7037 (n4048, n700, n_3630);
  not g7038 (n_3631, n4048);
  and g7039 (n4049, n704, n_3631);
  not g7040 (n_3632, n4049);
  and g7041 (n4050, n708, n_3632);
  not g7042 (n_3633, n4050);
  and g7043 (n4051, n712, n_3633);
  not g7044 (n_3634, n4051);
  and g7045 (n4052, n716, n_3634);
  not g7046 (n_3635, n4052);
  and g7047 (n4053, n720, n_3635);
  not g7048 (n_3636, n4053);
  and g7049 (n4054, n1484, n_3636);
  not g7050 (n_3637, n4054);
  and g7051 (n4055, n1486, n_3637);
  not g7052 (n_3638, n4055);
  and g7053 (n4056, n1750, n_3638);
  not g7054 (n_3639, n4056);
  and g7055 (n4057, n731, n_3639);
  not g7056 (n_3640, n4057);
  and g7057 (n4058, n735, n_3640);
  not g7058 (n_3641, n4058);
  and g7059 (n4059, n739, n_3641);
  not g7060 (n_3642, n4059);
  and g7061 (n4060, n743, n_3642);
  not g7062 (n_3643, n4060);
  and g7063 (n4061, n747, n_3643);
  not g7064 (n_3644, n4061);
  and g7065 (n4062, n751, n_3644);
  not g7066 (n_3645, n4062);
  and g7067 (n4063, n755, n_3645);
  not g7068 (n_3646, n4063);
  and g7069 (n4064, n759, n_3646);
  not g7070 (n_3647, n4064);
  and g7071 (n4065, n763, n_3647);
  not g7072 (n_3648, n4065);
  and g7073 (n4066, n767, n_3648);
  not g7074 (n_3649, n4066);
  and g7075 (n4067, n771, n_3649);
  not g7076 (n_3650, n4067);
  and g7077 (n4068, n775, n_3650);
  not g7078 (n_3651, n4068);
  and g7079 (n4069, n779, n_3651);
  not g7080 (n_3652, n4069);
  and g7081 (n4070, n783, n_3652);
  not g7082 (n_3653, n4070);
  and g7083 (n4071, n787, n_3653);
  not g7084 (n_3654, n4071);
  and g7085 (n4072, n791, n_3654);
  not g7086 (n_3655, n4072);
  and g7087 (n4073, n795, n_3655);
  not g7088 (n_3656, n4073);
  and g7089 (n4074, n799, n_3656);
  not g7090 (n_3657, n4074);
  and g7091 (n4075, n803, n_3657);
  and g7092 (n4076, \req[33] , n_659);
  not g7093 (n_3658, n4075);
  and g7094 (\grant[33] , n_3658, n4076);
  not g7095 (n_3659, n1147);
  and g7096 (n4078, n814, n_3659);
  not g7097 (n_3660, n4078);
  and g7098 (n4079, n819, n_3660);
  not g7099 (n_3661, n4079);
  and g7100 (n4080, n823, n_3661);
  not g7101 (n_3662, n4080);
  and g7102 (n4081, n827, n_3662);
  not g7103 (n_3663, n4081);
  and g7104 (n4082, n831, n_3663);
  not g7105 (n_3664, n4082);
  and g7106 (n4083, n835, n_3664);
  not g7107 (n_3665, n4083);
  and g7108 (n4084, n839, n_3665);
  not g7109 (n_3666, n4084);
  and g7110 (n4085, n843, n_3666);
  not g7111 (n_3667, n4085);
  and g7112 (n4086, n847, n_3667);
  not g7113 (n_3668, n4086);
  and g7114 (n4087, n851, n_3668);
  not g7115 (n_3669, n4087);
  and g7116 (n4088, n855, n_3669);
  not g7117 (n_3670, n4088);
  and g7118 (n4089, n859, n_3670);
  not g7119 (n_3671, n4089);
  and g7120 (n4090, n863, n_3671);
  not g7121 (n_3672, n4090);
  and g7122 (n4091, n867, n_3672);
  not g7123 (n_3673, n4091);
  and g7124 (n4092, n871, n_3673);
  not g7125 (n_3674, n4092);
  and g7126 (n4093, n875, n_3674);
  not g7127 (n_3675, n4093);
  and g7128 (n4094, n879, n_3675);
  not g7129 (n_3676, n4094);
  and g7130 (n4095, n883, n_3676);
  not g7131 (n_3677, n4095);
  and g7132 (n4096, n887, n_3677);
  not g7133 (n_3678, n4096);
  and g7134 (n4097, n891, n_3678);
  not g7135 (n_3679, n4097);
  and g7136 (n4098, n895, n_3679);
  not g7137 (n_3680, n4098);
  and g7138 (n4099, n899, n_3680);
  not g7139 (n_3681, n4099);
  and g7140 (n4100, n903, n_3681);
  not g7141 (n_3682, n4100);
  and g7142 (n4101, n907, n_3682);
  not g7143 (n_3683, n4101);
  and g7144 (n4102, n911, n_3683);
  not g7145 (n_3684, n4102);
  and g7146 (n4103, n915, n_3684);
  not g7147 (n_3685, n4103);
  and g7148 (n4104, n919, n_3685);
  not g7149 (n_3686, n4104);
  and g7150 (n4105, n923, n_3686);
  not g7151 (n_3687, n4105);
  and g7152 (n4106, n927, n_3687);
  not g7153 (n_3688, n4106);
  and g7154 (n4107, n931, n_3688);
  not g7155 (n_3689, n4107);
  and g7156 (n4108, n935, n_3689);
  not g7157 (n_3690, n4108);
  and g7158 (n4109, n939, n_3690);
  not g7159 (n_3691, n4109);
  and g7160 (n4110, n943, n_3691);
  not g7161 (n_3692, n4110);
  and g7162 (n4111, n947, n_3692);
  not g7163 (n_3693, n4111);
  and g7164 (n4112, n951, n_3693);
  not g7165 (n_3694, n4112);
  and g7166 (n4113, n955, n_3694);
  not g7167 (n_3695, n4113);
  and g7168 (n4114, n959, n_3695);
  not g7169 (n_3696, n4114);
  and g7170 (n4115, n963, n_3696);
  not g7171 (n_3697, n4115);
  and g7172 (n4116, n967, n_3697);
  not g7173 (n_3698, n4116);
  and g7174 (n4117, n971, n_3698);
  not g7175 (n_3699, n4117);
  and g7176 (n4118, n975, n_3699);
  not g7177 (n_3700, n4118);
  and g7178 (n4119, n979, n_3700);
  not g7179 (n_3701, n4119);
  and g7180 (n4120, n983, n_3701);
  not g7181 (n_3702, n4120);
  and g7182 (n4121, n987, n_3702);
  not g7183 (n_3703, n4121);
  and g7184 (n4122, n991, n_3703);
  not g7185 (n_3704, n4122);
  and g7186 (n4123, n995, n_3704);
  not g7187 (n_3705, n4123);
  and g7188 (n4124, n999, n_3705);
  not g7189 (n_3706, n4124);
  and g7190 (n4125, n1003, n_3706);
  not g7191 (n_3707, n4125);
  and g7192 (n4126, n1007, n_3707);
  not g7193 (n_3708, n4126);
  and g7194 (n4127, n1011, n_3708);
  not g7195 (n_3709, n4127);
  and g7196 (n4128, n1015, n_3709);
  not g7197 (n_3710, n4128);
  and g7198 (n4129, n1019, n_3710);
  not g7199 (n_3711, n4129);
  and g7200 (n4130, n1023, n_3711);
  not g7201 (n_3712, n4130);
  and g7202 (n4131, n1027, n_3712);
  not g7203 (n_3713, n4131);
  and g7204 (n4132, n1031, n_3713);
  not g7205 (n_3714, n4132);
  and g7206 (n4133, n1035, n_3714);
  not g7207 (n_3715, n4133);
  and g7208 (n4134, n1039, n_3715);
  not g7209 (n_3716, n4134);
  and g7210 (n4135, n1043, n_3716);
  not g7211 (n_3717, n4135);
  and g7212 (n4136, n1047, n_3717);
  not g7213 (n_3718, n4136);
  and g7214 (n4137, n1051, n_3718);
  not g7215 (n_3719, n4137);
  and g7216 (n4138, n1055, n_3719);
  not g7217 (n_3720, n4138);
  and g7218 (n4139, n1059, n_3720);
  not g7219 (n_3721, n4139);
  and g7220 (n4140, n1574, n_3721);
  not g7221 (n_3722, n4140);
  and g7222 (n4141, n1576, n_3722);
  not g7223 (n_3723, n4141);
  and g7224 (n4142, n1837, n_3723);
  not g7225 (n_3724, n4142);
  and g7226 (n4143, n1068, n_3724);
  not g7227 (n_3725, n4143);
  and g7228 (n4144, n1072, n_3725);
  not g7229 (n_3726, n4144);
  and g7230 (n4145, n1076, n_3726);
  not g7231 (n_3727, n4145);
  and g7232 (n4146, n1080, n_3727);
  not g7233 (n_3728, n4146);
  and g7234 (n4147, n1084, n_3728);
  not g7235 (n_3729, n4147);
  and g7236 (n4148, n1088, n_3729);
  not g7237 (n_3730, n4148);
  and g7238 (n4149, n1092, n_3730);
  not g7239 (n_3731, n4149);
  and g7240 (n4150, n1096, n_3731);
  not g7241 (n_3732, n4150);
  and g7242 (n4151, n1100, n_3732);
  not g7243 (n_3733, n4151);
  and g7244 (n4152, n1104, n_3733);
  not g7245 (n_3734, n4152);
  and g7246 (n4153, n1108, n_3734);
  not g7247 (n_3735, n4153);
  and g7248 (n4154, n1112, n_3735);
  not g7249 (n_3736, n4154);
  and g7250 (n4155, n1116, n_3736);
  not g7251 (n_3737, n4155);
  and g7252 (n4156, n1120, n_3737);
  not g7253 (n_3738, n4156);
  and g7254 (n4157, n1124, n_3738);
  not g7255 (n_3739, n4157);
  and g7256 (n4158, n1128, n_3739);
  not g7257 (n_3740, n4158);
  and g7258 (n4159, n1132, n_3740);
  not g7259 (n_3741, n4159);
  and g7260 (n4160, n1136, n_3741);
  not g7261 (n_3742, n4160);
  and g7262 (n4161, n1140, n_3742);
  and g7263 (n4162, \req[34] , n_891);
  not g7264 (n_3743, n4161);
  and g7265 (\grant[34] , n_3743, n4162);
  not g7266 (n_3744, n479);
  and g7267 (n4164, n_3744, n1151);
  not g7268 (n_3745, n4164);
  and g7269 (n4165, n1156, n_3745);
  not g7270 (n_3746, n4165);
  and g7271 (n4166, n1160, n_3746);
  not g7272 (n_3747, n4166);
  and g7273 (n4167, n1164, n_3747);
  not g7274 (n_3748, n4167);
  and g7275 (n4168, n1168, n_3748);
  not g7276 (n_3749, n4168);
  and g7277 (n4169, n1172, n_3749);
  not g7278 (n_3750, n4169);
  and g7279 (n4170, n1176, n_3750);
  not g7280 (n_3751, n4170);
  and g7281 (n4171, n1180, n_3751);
  not g7282 (n_3752, n4171);
  and g7283 (n4172, n1184, n_3752);
  not g7284 (n_3753, n4172);
  and g7285 (n4173, n1188, n_3753);
  not g7286 (n_3754, n4173);
  and g7287 (n4174, n1192, n_3754);
  not g7288 (n_3755, n4174);
  and g7289 (n4175, n1196, n_3755);
  not g7290 (n_3756, n4175);
  and g7291 (n4176, n1200, n_3756);
  not g7292 (n_3757, n4176);
  and g7293 (n4177, n1204, n_3757);
  not g7294 (n_3758, n4177);
  and g7295 (n4178, n1208, n_3758);
  not g7296 (n_3759, n4178);
  and g7297 (n4179, n1212, n_3759);
  not g7298 (n_3760, n4179);
  and g7299 (n4180, n1216, n_3760);
  not g7300 (n_3761, n4180);
  and g7301 (n4181, n1220, n_3761);
  not g7302 (n_3762, n4181);
  and g7303 (n4182, n1224, n_3762);
  not g7304 (n_3763, n4182);
  and g7305 (n4183, n1228, n_3763);
  not g7306 (n_3764, n4183);
  and g7307 (n4184, n1232, n_3764);
  not g7308 (n_3765, n4184);
  and g7309 (n4185, n1236, n_3765);
  not g7310 (n_3766, n4185);
  and g7311 (n4186, n1240, n_3766);
  not g7312 (n_3767, n4186);
  and g7313 (n4187, n1244, n_3767);
  not g7314 (n_3768, n4187);
  and g7315 (n4188, n1248, n_3768);
  not g7316 (n_3769, n4188);
  and g7317 (n4189, n1252, n_3769);
  not g7318 (n_3770, n4189);
  and g7319 (n4190, n1256, n_3770);
  not g7320 (n_3771, n4190);
  and g7321 (n4191, n1260, n_3771);
  not g7322 (n_3772, n4191);
  and g7323 (n4192, n1264, n_3772);
  not g7324 (n_3773, n4192);
  and g7325 (n4193, n1268, n_3773);
  not g7326 (n_3774, n4193);
  and g7327 (n4194, n1272, n_3774);
  not g7328 (n_3775, n4194);
  and g7329 (n4195, n1276, n_3775);
  not g7330 (n_3776, n4195);
  and g7331 (n4196, n1280, n_3776);
  not g7332 (n_3777, n4196);
  and g7333 (n4197, n1284, n_3777);
  not g7334 (n_3778, n4197);
  and g7335 (n4198, n1288, n_3778);
  not g7336 (n_3779, n4198);
  and g7337 (n4199, n1292, n_3779);
  not g7338 (n_3780, n4199);
  and g7339 (n4200, n1296, n_3780);
  not g7340 (n_3781, n4200);
  and g7341 (n4201, n1300, n_3781);
  not g7342 (n_3782, n4201);
  and g7343 (n4202, n1304, n_3782);
  not g7344 (n_3783, n4202);
  and g7345 (n4203, n1308, n_3783);
  not g7346 (n_3784, n4203);
  and g7347 (n4204, n1312, n_3784);
  not g7348 (n_3785, n4204);
  and g7349 (n4205, n1316, n_3785);
  not g7350 (n_3786, n4205);
  and g7351 (n4206, n1320, n_3786);
  not g7352 (n_3787, n4206);
  and g7353 (n4207, n1324, n_3787);
  not g7354 (n_3788, n4207);
  and g7355 (n4208, n1328, n_3788);
  not g7356 (n_3789, n4208);
  and g7357 (n4209, n1332, n_3789);
  not g7358 (n_3790, n4209);
  and g7359 (n4210, n1336, n_3790);
  not g7360 (n_3791, n4210);
  and g7361 (n4211, n1340, n_3791);
  not g7362 (n_3792, n4211);
  and g7363 (n4212, n1344, n_3792);
  not g7364 (n_3793, n4212);
  and g7365 (n4213, n1348, n_3793);
  not g7366 (n_3794, n4213);
  and g7367 (n4214, n1352, n_3794);
  not g7368 (n_3795, n4214);
  and g7369 (n4215, n1356, n_3795);
  not g7370 (n_3796, n4215);
  and g7371 (n4216, n1360, n_3796);
  not g7372 (n_3797, n4216);
  and g7373 (n4217, n1364, n_3797);
  not g7374 (n_3798, n4217);
  and g7375 (n4218, n1368, n_3798);
  not g7376 (n_3799, n4218);
  and g7377 (n4219, n1372, n_3799);
  not g7378 (n_3800, n4219);
  and g7379 (n4220, n1376, n_3800);
  not g7380 (n_3801, n4220);
  and g7381 (n4221, n1380, n_3801);
  not g7382 (n_3802, n4221);
  and g7383 (n4222, n1384, n_3802);
  not g7384 (n_3803, n4222);
  and g7385 (n4223, n1388, n_3803);
  not g7386 (n_3804, n4223);
  and g7387 (n4224, n1392, n_3804);
  not g7388 (n_3805, n4224);
  and g7389 (n4225, n1396, n_3805);
  not g7390 (n_3806, n4225);
  and g7391 (n4226, n1663, n_3806);
  not g7392 (n_3807, n4226);
  and g7393 (n4227, n392, n_3807);
  not g7394 (n_3808, n4227);
  and g7395 (n4228, n396, n_3808);
  not g7396 (n_3809, n4228);
  and g7397 (n4229, n400, n_3809);
  not g7398 (n_3810, n4229);
  and g7399 (n4230, n404, n_3810);
  not g7400 (n_3811, n4230);
  and g7401 (n4231, n408, n_3811);
  not g7402 (n_3812, n4231);
  and g7403 (n4232, n412, n_3812);
  not g7404 (n_3813, n4232);
  and g7405 (n4233, n416, n_3813);
  not g7406 (n_3814, n4233);
  and g7407 (n4234, n420, n_3814);
  not g7408 (n_3815, n4234);
  and g7409 (n4235, n424, n_3815);
  not g7410 (n_3816, n4235);
  and g7411 (n4236, n428, n_3816);
  not g7412 (n_3817, n4236);
  and g7413 (n4237, n432, n_3817);
  not g7414 (n_3818, n4237);
  and g7415 (n4238, n436, n_3818);
  not g7416 (n_3819, n4238);
  and g7417 (n4239, n440, n_3819);
  not g7418 (n_3820, n4239);
  and g7419 (n4240, n444, n_3820);
  not g7420 (n_3821, n4240);
  and g7421 (n4241, n448, n_3821);
  not g7422 (n_3822, n4241);
  and g7423 (n4242, n452, n_3822);
  not g7424 (n_3823, n4242);
  and g7425 (n4243, n456, n_3823);
  not g7426 (n_3824, n4243);
  and g7427 (n4244, n460, n_3824);
  not g7428 (n_3825, n4244);
  and g7429 (n4245, n464, n_3825);
  not g7430 (n_3826, n4245);
  and g7431 (n4246, n468, n_3826);
  not g7432 (n_3827, n4246);
  and g7433 (n4247, n472, n_3827);
  and g7434 (n4248, \req[35] , n_164);
  not g7435 (n_3828, n4247);
  and g7436 (\grant[35] , n_3828, n4248);
  not g7437 (n_3829, n818);
  and g7438 (n4250, n483, n_3829);
  not g7439 (n_3830, n4250);
  and g7440 (n4251, n488, n_3830);
  not g7441 (n_3831, n4251);
  and g7442 (n4252, n492, n_3831);
  not g7443 (n_3832, n4252);
  and g7444 (n4253, n496, n_3832);
  not g7445 (n_3833, n4253);
  and g7446 (n4254, n500, n_3833);
  not g7447 (n_3834, n4254);
  and g7448 (n4255, n504, n_3834);
  not g7449 (n_3835, n4255);
  and g7450 (n4256, n508, n_3835);
  not g7451 (n_3836, n4256);
  and g7452 (n4257, n512, n_3836);
  not g7453 (n_3837, n4257);
  and g7454 (n4258, n516, n_3837);
  not g7455 (n_3838, n4258);
  and g7456 (n4259, n520, n_3838);
  not g7457 (n_3839, n4259);
  and g7458 (n4260, n524, n_3839);
  not g7459 (n_3840, n4260);
  and g7460 (n4261, n528, n_3840);
  not g7461 (n_3841, n4261);
  and g7462 (n4262, n532, n_3841);
  not g7463 (n_3842, n4262);
  and g7464 (n4263, n536, n_3842);
  not g7465 (n_3843, n4263);
  and g7466 (n4264, n540, n_3843);
  not g7467 (n_3844, n4264);
  and g7468 (n4265, n544, n_3844);
  not g7469 (n_3845, n4265);
  and g7470 (n4266, n548, n_3845);
  not g7471 (n_3846, n4266);
  and g7472 (n4267, n552, n_3846);
  not g7473 (n_3847, n4267);
  and g7474 (n4268, n556, n_3847);
  not g7475 (n_3848, n4268);
  and g7476 (n4269, n560, n_3848);
  not g7477 (n_3849, n4269);
  and g7478 (n4270, n564, n_3849);
  not g7479 (n_3850, n4270);
  and g7480 (n4271, n568, n_3850);
  not g7481 (n_3851, n4271);
  and g7482 (n4272, n572, n_3851);
  not g7483 (n_3852, n4272);
  and g7484 (n4273, n576, n_3852);
  not g7485 (n_3853, n4273);
  and g7486 (n4274, n580, n_3853);
  not g7487 (n_3854, n4274);
  and g7488 (n4275, n584, n_3854);
  not g7489 (n_3855, n4275);
  and g7490 (n4276, n588, n_3855);
  not g7491 (n_3856, n4276);
  and g7492 (n4277, n592, n_3856);
  not g7493 (n_3857, n4277);
  and g7494 (n4278, n596, n_3857);
  not g7495 (n_3858, n4278);
  and g7496 (n4279, n600, n_3858);
  not g7497 (n_3859, n4279);
  and g7498 (n4280, n604, n_3859);
  not g7499 (n_3860, n4280);
  and g7500 (n4281, n608, n_3860);
  not g7501 (n_3861, n4281);
  and g7502 (n4282, n612, n_3861);
  not g7503 (n_3862, n4282);
  and g7504 (n4283, n616, n_3862);
  not g7505 (n_3863, n4283);
  and g7506 (n4284, n620, n_3863);
  not g7507 (n_3864, n4284);
  and g7508 (n4285, n624, n_3864);
  not g7509 (n_3865, n4285);
  and g7510 (n4286, n628, n_3865);
  not g7511 (n_3866, n4286);
  and g7512 (n4287, n632, n_3866);
  not g7513 (n_3867, n4287);
  and g7514 (n4288, n636, n_3867);
  not g7515 (n_3868, n4288);
  and g7516 (n4289, n640, n_3868);
  not g7517 (n_3869, n4289);
  and g7518 (n4290, n644, n_3869);
  not g7519 (n_3870, n4290);
  and g7520 (n4291, n648, n_3870);
  not g7521 (n_3871, n4291);
  and g7522 (n4292, n652, n_3871);
  not g7523 (n_3872, n4292);
  and g7524 (n4293, n656, n_3872);
  not g7525 (n_3873, n4293);
  and g7526 (n4294, n660, n_3873);
  not g7527 (n_3874, n4294);
  and g7528 (n4295, n664, n_3874);
  not g7529 (n_3875, n4295);
  and g7530 (n4296, n668, n_3875);
  not g7531 (n_3876, n4296);
  and g7532 (n4297, n672, n_3876);
  not g7533 (n_3877, n4297);
  and g7534 (n4298, n676, n_3877);
  not g7535 (n_3878, n4298);
  and g7536 (n4299, n680, n_3878);
  not g7537 (n_3879, n4299);
  and g7538 (n4300, n684, n_3879);
  not g7539 (n_3880, n4300);
  and g7540 (n4301, n688, n_3880);
  not g7541 (n_3881, n4301);
  and g7542 (n4302, n692, n_3881);
  not g7543 (n_3882, n4302);
  and g7544 (n4303, n696, n_3882);
  not g7545 (n_3883, n4303);
  and g7546 (n4304, n700, n_3883);
  not g7547 (n_3884, n4304);
  and g7548 (n4305, n704, n_3884);
  not g7549 (n_3885, n4305);
  and g7550 (n4306, n708, n_3885);
  not g7551 (n_3886, n4306);
  and g7552 (n4307, n712, n_3886);
  not g7553 (n_3887, n4307);
  and g7554 (n4308, n716, n_3887);
  not g7555 (n_3888, n4308);
  and g7556 (n4309, n720, n_3888);
  not g7557 (n_3889, n4309);
  and g7558 (n4310, n1484, n_3889);
  not g7559 (n_3890, n4310);
  and g7560 (n4311, n1486, n_3890);
  not g7561 (n_3891, n4311);
  and g7562 (n4312, n1750, n_3891);
  not g7563 (n_3892, n4312);
  and g7564 (n4313, n731, n_3892);
  not g7565 (n_3893, n4313);
  and g7566 (n4314, n735, n_3893);
  not g7567 (n_3894, n4314);
  and g7568 (n4315, n739, n_3894);
  not g7569 (n_3895, n4315);
  and g7570 (n4316, n743, n_3895);
  not g7571 (n_3896, n4316);
  and g7572 (n4317, n747, n_3896);
  not g7573 (n_3897, n4317);
  and g7574 (n4318, n751, n_3897);
  not g7575 (n_3898, n4318);
  and g7576 (n4319, n755, n_3898);
  not g7577 (n_3899, n4319);
  and g7578 (n4320, n759, n_3899);
  not g7579 (n_3900, n4320);
  and g7580 (n4321, n763, n_3900);
  not g7581 (n_3901, n4321);
  and g7582 (n4322, n767, n_3901);
  not g7583 (n_3902, n4322);
  and g7584 (n4323, n771, n_3902);
  not g7585 (n_3903, n4323);
  and g7586 (n4324, n775, n_3903);
  not g7587 (n_3904, n4324);
  and g7588 (n4325, n779, n_3904);
  not g7589 (n_3905, n4325);
  and g7590 (n4326, n783, n_3905);
  not g7591 (n_3906, n4326);
  and g7592 (n4327, n787, n_3906);
  not g7593 (n_3907, n4327);
  and g7594 (n4328, n791, n_3907);
  not g7595 (n_3908, n4328);
  and g7596 (n4329, n795, n_3908);
  not g7597 (n_3909, n4329);
  and g7598 (n4330, n799, n_3909);
  not g7599 (n_3910, n4330);
  and g7600 (n4331, n803, n_3910);
  not g7601 (n_3911, n4331);
  and g7602 (n4332, n807, n_3911);
  not g7603 (n_3912, n4332);
  and g7604 (n4333, n811, n_3912);
  and g7605 (n4334, \req[36] , n_665);
  not g7606 (n_3913, n4333);
  and g7607 (\grant[36] , n_3913, n4334);
  not g7608 (n_3914, n1155);
  and g7609 (n4336, n822, n_3914);
  not g7610 (n_3915, n4336);
  and g7611 (n4337, n827, n_3915);
  not g7612 (n_3916, n4337);
  and g7613 (n4338, n831, n_3916);
  not g7614 (n_3917, n4338);
  and g7615 (n4339, n835, n_3917);
  not g7616 (n_3918, n4339);
  and g7617 (n4340, n839, n_3918);
  not g7618 (n_3919, n4340);
  and g7619 (n4341, n843, n_3919);
  not g7620 (n_3920, n4341);
  and g7621 (n4342, n847, n_3920);
  not g7622 (n_3921, n4342);
  and g7623 (n4343, n851, n_3921);
  not g7624 (n_3922, n4343);
  and g7625 (n4344, n855, n_3922);
  not g7626 (n_3923, n4344);
  and g7627 (n4345, n859, n_3923);
  not g7628 (n_3924, n4345);
  and g7629 (n4346, n863, n_3924);
  not g7630 (n_3925, n4346);
  and g7631 (n4347, n867, n_3925);
  not g7632 (n_3926, n4347);
  and g7633 (n4348, n871, n_3926);
  not g7634 (n_3927, n4348);
  and g7635 (n4349, n875, n_3927);
  not g7636 (n_3928, n4349);
  and g7637 (n4350, n879, n_3928);
  not g7638 (n_3929, n4350);
  and g7639 (n4351, n883, n_3929);
  not g7640 (n_3930, n4351);
  and g7641 (n4352, n887, n_3930);
  not g7642 (n_3931, n4352);
  and g7643 (n4353, n891, n_3931);
  not g7644 (n_3932, n4353);
  and g7645 (n4354, n895, n_3932);
  not g7646 (n_3933, n4354);
  and g7647 (n4355, n899, n_3933);
  not g7648 (n_3934, n4355);
  and g7649 (n4356, n903, n_3934);
  not g7650 (n_3935, n4356);
  and g7651 (n4357, n907, n_3935);
  not g7652 (n_3936, n4357);
  and g7653 (n4358, n911, n_3936);
  not g7654 (n_3937, n4358);
  and g7655 (n4359, n915, n_3937);
  not g7656 (n_3938, n4359);
  and g7657 (n4360, n919, n_3938);
  not g7658 (n_3939, n4360);
  and g7659 (n4361, n923, n_3939);
  not g7660 (n_3940, n4361);
  and g7661 (n4362, n927, n_3940);
  not g7662 (n_3941, n4362);
  and g7663 (n4363, n931, n_3941);
  not g7664 (n_3942, n4363);
  and g7665 (n4364, n935, n_3942);
  not g7666 (n_3943, n4364);
  and g7667 (n4365, n939, n_3943);
  not g7668 (n_3944, n4365);
  and g7669 (n4366, n943, n_3944);
  not g7670 (n_3945, n4366);
  and g7671 (n4367, n947, n_3945);
  not g7672 (n_3946, n4367);
  and g7673 (n4368, n951, n_3946);
  not g7674 (n_3947, n4368);
  and g7675 (n4369, n955, n_3947);
  not g7676 (n_3948, n4369);
  and g7677 (n4370, n959, n_3948);
  not g7678 (n_3949, n4370);
  and g7679 (n4371, n963, n_3949);
  not g7680 (n_3950, n4371);
  and g7681 (n4372, n967, n_3950);
  not g7682 (n_3951, n4372);
  and g7683 (n4373, n971, n_3951);
  not g7684 (n_3952, n4373);
  and g7685 (n4374, n975, n_3952);
  not g7686 (n_3953, n4374);
  and g7687 (n4375, n979, n_3953);
  not g7688 (n_3954, n4375);
  and g7689 (n4376, n983, n_3954);
  not g7690 (n_3955, n4376);
  and g7691 (n4377, n987, n_3955);
  not g7692 (n_3956, n4377);
  and g7693 (n4378, n991, n_3956);
  not g7694 (n_3957, n4378);
  and g7695 (n4379, n995, n_3957);
  not g7696 (n_3958, n4379);
  and g7697 (n4380, n999, n_3958);
  not g7698 (n_3959, n4380);
  and g7699 (n4381, n1003, n_3959);
  not g7700 (n_3960, n4381);
  and g7701 (n4382, n1007, n_3960);
  not g7702 (n_3961, n4382);
  and g7703 (n4383, n1011, n_3961);
  not g7704 (n_3962, n4383);
  and g7705 (n4384, n1015, n_3962);
  not g7706 (n_3963, n4384);
  and g7707 (n4385, n1019, n_3963);
  not g7708 (n_3964, n4385);
  and g7709 (n4386, n1023, n_3964);
  not g7710 (n_3965, n4386);
  and g7711 (n4387, n1027, n_3965);
  not g7712 (n_3966, n4387);
  and g7713 (n4388, n1031, n_3966);
  not g7714 (n_3967, n4388);
  and g7715 (n4389, n1035, n_3967);
  not g7716 (n_3968, n4389);
  and g7717 (n4390, n1039, n_3968);
  not g7718 (n_3969, n4390);
  and g7719 (n4391, n1043, n_3969);
  not g7720 (n_3970, n4391);
  and g7721 (n4392, n1047, n_3970);
  not g7722 (n_3971, n4392);
  and g7723 (n4393, n1051, n_3971);
  not g7724 (n_3972, n4393);
  and g7725 (n4394, n1055, n_3972);
  not g7726 (n_3973, n4394);
  and g7727 (n4395, n1059, n_3973);
  not g7728 (n_3974, n4395);
  and g7729 (n4396, n1574, n_3974);
  not g7730 (n_3975, n4396);
  and g7731 (n4397, n1576, n_3975);
  not g7732 (n_3976, n4397);
  and g7733 (n4398, n1837, n_3976);
  not g7734 (n_3977, n4398);
  and g7735 (n4399, n1068, n_3977);
  not g7736 (n_3978, n4399);
  and g7737 (n4400, n1072, n_3978);
  not g7738 (n_3979, n4400);
  and g7739 (n4401, n1076, n_3979);
  not g7740 (n_3980, n4401);
  and g7741 (n4402, n1080, n_3980);
  not g7742 (n_3981, n4402);
  and g7743 (n4403, n1084, n_3981);
  not g7744 (n_3982, n4403);
  and g7745 (n4404, n1088, n_3982);
  not g7746 (n_3983, n4404);
  and g7747 (n4405, n1092, n_3983);
  not g7748 (n_3984, n4405);
  and g7749 (n4406, n1096, n_3984);
  not g7750 (n_3985, n4406);
  and g7751 (n4407, n1100, n_3985);
  not g7752 (n_3986, n4407);
  and g7753 (n4408, n1104, n_3986);
  not g7754 (n_3987, n4408);
  and g7755 (n4409, n1108, n_3987);
  not g7756 (n_3988, n4409);
  and g7757 (n4410, n1112, n_3988);
  not g7758 (n_3989, n4410);
  and g7759 (n4411, n1116, n_3989);
  not g7760 (n_3990, n4411);
  and g7761 (n4412, n1120, n_3990);
  not g7762 (n_3991, n4412);
  and g7763 (n4413, n1124, n_3991);
  not g7764 (n_3992, n4413);
  and g7765 (n4414, n1128, n_3992);
  not g7766 (n_3993, n4414);
  and g7767 (n4415, n1132, n_3993);
  not g7768 (n_3994, n4415);
  and g7769 (n4416, n1136, n_3994);
  not g7770 (n_3995, n4416);
  and g7771 (n4417, n1140, n_3995);
  not g7772 (n_3996, n4417);
  and g7773 (n4418, n1144, n_3996);
  not g7774 (n_3997, n4418);
  and g7775 (n4419, n1148, n_3997);
  and g7776 (n4420, \req[37] , n_895);
  not g7777 (n_3998, n4419);
  and g7778 (\grant[37] , n_3998, n4420);
  not g7779 (n_3999, n487);
  and g7780 (n4422, n_3999, n1159);
  not g7781 (n_4000, n4422);
  and g7782 (n4423, n1164, n_4000);
  not g7783 (n_4001, n4423);
  and g7784 (n4424, n1168, n_4001);
  not g7785 (n_4002, n4424);
  and g7786 (n4425, n1172, n_4002);
  not g7787 (n_4003, n4425);
  and g7788 (n4426, n1176, n_4003);
  not g7789 (n_4004, n4426);
  and g7790 (n4427, n1180, n_4004);
  not g7791 (n_4005, n4427);
  and g7792 (n4428, n1184, n_4005);
  not g7793 (n_4006, n4428);
  and g7794 (n4429, n1188, n_4006);
  not g7795 (n_4007, n4429);
  and g7796 (n4430, n1192, n_4007);
  not g7797 (n_4008, n4430);
  and g7798 (n4431, n1196, n_4008);
  not g7799 (n_4009, n4431);
  and g7800 (n4432, n1200, n_4009);
  not g7801 (n_4010, n4432);
  and g7802 (n4433, n1204, n_4010);
  not g7803 (n_4011, n4433);
  and g7804 (n4434, n1208, n_4011);
  not g7805 (n_4012, n4434);
  and g7806 (n4435, n1212, n_4012);
  not g7807 (n_4013, n4435);
  and g7808 (n4436, n1216, n_4013);
  not g7809 (n_4014, n4436);
  and g7810 (n4437, n1220, n_4014);
  not g7811 (n_4015, n4437);
  and g7812 (n4438, n1224, n_4015);
  not g7813 (n_4016, n4438);
  and g7814 (n4439, n1228, n_4016);
  not g7815 (n_4017, n4439);
  and g7816 (n4440, n1232, n_4017);
  not g7817 (n_4018, n4440);
  and g7818 (n4441, n1236, n_4018);
  not g7819 (n_4019, n4441);
  and g7820 (n4442, n1240, n_4019);
  not g7821 (n_4020, n4442);
  and g7822 (n4443, n1244, n_4020);
  not g7823 (n_4021, n4443);
  and g7824 (n4444, n1248, n_4021);
  not g7825 (n_4022, n4444);
  and g7826 (n4445, n1252, n_4022);
  not g7827 (n_4023, n4445);
  and g7828 (n4446, n1256, n_4023);
  not g7829 (n_4024, n4446);
  and g7830 (n4447, n1260, n_4024);
  not g7831 (n_4025, n4447);
  and g7832 (n4448, n1264, n_4025);
  not g7833 (n_4026, n4448);
  and g7834 (n4449, n1268, n_4026);
  not g7835 (n_4027, n4449);
  and g7836 (n4450, n1272, n_4027);
  not g7837 (n_4028, n4450);
  and g7838 (n4451, n1276, n_4028);
  not g7839 (n_4029, n4451);
  and g7840 (n4452, n1280, n_4029);
  not g7841 (n_4030, n4452);
  and g7842 (n4453, n1284, n_4030);
  not g7843 (n_4031, n4453);
  and g7844 (n4454, n1288, n_4031);
  not g7845 (n_4032, n4454);
  and g7846 (n4455, n1292, n_4032);
  not g7847 (n_4033, n4455);
  and g7848 (n4456, n1296, n_4033);
  not g7849 (n_4034, n4456);
  and g7850 (n4457, n1300, n_4034);
  not g7851 (n_4035, n4457);
  and g7852 (n4458, n1304, n_4035);
  not g7853 (n_4036, n4458);
  and g7854 (n4459, n1308, n_4036);
  not g7855 (n_4037, n4459);
  and g7856 (n4460, n1312, n_4037);
  not g7857 (n_4038, n4460);
  and g7858 (n4461, n1316, n_4038);
  not g7859 (n_4039, n4461);
  and g7860 (n4462, n1320, n_4039);
  not g7861 (n_4040, n4462);
  and g7862 (n4463, n1324, n_4040);
  not g7863 (n_4041, n4463);
  and g7864 (n4464, n1328, n_4041);
  not g7865 (n_4042, n4464);
  and g7866 (n4465, n1332, n_4042);
  not g7867 (n_4043, n4465);
  and g7868 (n4466, n1336, n_4043);
  not g7869 (n_4044, n4466);
  and g7870 (n4467, n1340, n_4044);
  not g7871 (n_4045, n4467);
  and g7872 (n4468, n1344, n_4045);
  not g7873 (n_4046, n4468);
  and g7874 (n4469, n1348, n_4046);
  not g7875 (n_4047, n4469);
  and g7876 (n4470, n1352, n_4047);
  not g7877 (n_4048, n4470);
  and g7878 (n4471, n1356, n_4048);
  not g7879 (n_4049, n4471);
  and g7880 (n4472, n1360, n_4049);
  not g7881 (n_4050, n4472);
  and g7882 (n4473, n1364, n_4050);
  not g7883 (n_4051, n4473);
  and g7884 (n4474, n1368, n_4051);
  not g7885 (n_4052, n4474);
  and g7886 (n4475, n1372, n_4052);
  not g7887 (n_4053, n4475);
  and g7888 (n4476, n1376, n_4053);
  not g7889 (n_4054, n4476);
  and g7890 (n4477, n1380, n_4054);
  not g7891 (n_4055, n4477);
  and g7892 (n4478, n1384, n_4055);
  not g7893 (n_4056, n4478);
  and g7894 (n4479, n1388, n_4056);
  not g7895 (n_4057, n4479);
  and g7896 (n4480, n1392, n_4057);
  not g7897 (n_4058, n4480);
  and g7898 (n4481, n1396, n_4058);
  not g7899 (n_4059, n4481);
  and g7900 (n4482, n1663, n_4059);
  not g7901 (n_4060, n4482);
  and g7902 (n4483, n392, n_4060);
  not g7903 (n_4061, n4483);
  and g7904 (n4484, n396, n_4061);
  not g7905 (n_4062, n4484);
  and g7906 (n4485, n400, n_4062);
  not g7907 (n_4063, n4485);
  and g7908 (n4486, n404, n_4063);
  not g7909 (n_4064, n4486);
  and g7910 (n4487, n408, n_4064);
  not g7911 (n_4065, n4487);
  and g7912 (n4488, n412, n_4065);
  not g7913 (n_4066, n4488);
  and g7914 (n4489, n416, n_4066);
  not g7915 (n_4067, n4489);
  and g7916 (n4490, n420, n_4067);
  not g7917 (n_4068, n4490);
  and g7918 (n4491, n424, n_4068);
  not g7919 (n_4069, n4491);
  and g7920 (n4492, n428, n_4069);
  not g7921 (n_4070, n4492);
  and g7922 (n4493, n432, n_4070);
  not g7923 (n_4071, n4493);
  and g7924 (n4494, n436, n_4071);
  not g7925 (n_4072, n4494);
  and g7926 (n4495, n440, n_4072);
  not g7927 (n_4073, n4495);
  and g7928 (n4496, n444, n_4073);
  not g7929 (n_4074, n4496);
  and g7930 (n4497, n448, n_4074);
  not g7931 (n_4075, n4497);
  and g7932 (n4498, n452, n_4075);
  not g7933 (n_4076, n4498);
  and g7934 (n4499, n456, n_4076);
  not g7935 (n_4077, n4499);
  and g7936 (n4500, n460, n_4077);
  not g7937 (n_4078, n4500);
  and g7938 (n4501, n464, n_4078);
  not g7939 (n_4079, n4501);
  and g7940 (n4502, n468, n_4079);
  not g7941 (n_4080, n4502);
  and g7942 (n4503, n472, n_4080);
  not g7943 (n_4081, n4503);
  and g7944 (n4504, n476, n_4081);
  not g7945 (n_4082, n4504);
  and g7946 (n4505, n480, n_4082);
  and g7947 (n4506, \req[38] , n_178);
  not g7948 (n_4083, n4505);
  and g7949 (\grant[38] , n_4083, n4506);
  not g7950 (n_4084, n826);
  and g7951 (n4508, n491, n_4084);
  not g7952 (n_4085, n4508);
  and g7953 (n4509, n496, n_4085);
  not g7954 (n_4086, n4509);
  and g7955 (n4510, n500, n_4086);
  not g7956 (n_4087, n4510);
  and g7957 (n4511, n504, n_4087);
  not g7958 (n_4088, n4511);
  and g7959 (n4512, n508, n_4088);
  not g7960 (n_4089, n4512);
  and g7961 (n4513, n512, n_4089);
  not g7962 (n_4090, n4513);
  and g7963 (n4514, n516, n_4090);
  not g7964 (n_4091, n4514);
  and g7965 (n4515, n520, n_4091);
  not g7966 (n_4092, n4515);
  and g7967 (n4516, n524, n_4092);
  not g7968 (n_4093, n4516);
  and g7969 (n4517, n528, n_4093);
  not g7970 (n_4094, n4517);
  and g7971 (n4518, n532, n_4094);
  not g7972 (n_4095, n4518);
  and g7973 (n4519, n536, n_4095);
  not g7974 (n_4096, n4519);
  and g7975 (n4520, n540, n_4096);
  not g7976 (n_4097, n4520);
  and g7977 (n4521, n544, n_4097);
  not g7978 (n_4098, n4521);
  and g7979 (n4522, n548, n_4098);
  not g7980 (n_4099, n4522);
  and g7981 (n4523, n552, n_4099);
  not g7982 (n_4100, n4523);
  and g7983 (n4524, n556, n_4100);
  not g7984 (n_4101, n4524);
  and g7985 (n4525, n560, n_4101);
  not g7986 (n_4102, n4525);
  and g7987 (n4526, n564, n_4102);
  not g7988 (n_4103, n4526);
  and g7989 (n4527, n568, n_4103);
  not g7990 (n_4104, n4527);
  and g7991 (n4528, n572, n_4104);
  not g7992 (n_4105, n4528);
  and g7993 (n4529, n576, n_4105);
  not g7994 (n_4106, n4529);
  and g7995 (n4530, n580, n_4106);
  not g7996 (n_4107, n4530);
  and g7997 (n4531, n584, n_4107);
  not g7998 (n_4108, n4531);
  and g7999 (n4532, n588, n_4108);
  not g8000 (n_4109, n4532);
  and g8001 (n4533, n592, n_4109);
  not g8002 (n_4110, n4533);
  and g8003 (n4534, n596, n_4110);
  not g8004 (n_4111, n4534);
  and g8005 (n4535, n600, n_4111);
  not g8006 (n_4112, n4535);
  and g8007 (n4536, n604, n_4112);
  not g8008 (n_4113, n4536);
  and g8009 (n4537, n608, n_4113);
  not g8010 (n_4114, n4537);
  and g8011 (n4538, n612, n_4114);
  not g8012 (n_4115, n4538);
  and g8013 (n4539, n616, n_4115);
  not g8014 (n_4116, n4539);
  and g8015 (n4540, n620, n_4116);
  not g8016 (n_4117, n4540);
  and g8017 (n4541, n624, n_4117);
  not g8018 (n_4118, n4541);
  and g8019 (n4542, n628, n_4118);
  not g8020 (n_4119, n4542);
  and g8021 (n4543, n632, n_4119);
  not g8022 (n_4120, n4543);
  and g8023 (n4544, n636, n_4120);
  not g8024 (n_4121, n4544);
  and g8025 (n4545, n640, n_4121);
  not g8026 (n_4122, n4545);
  and g8027 (n4546, n644, n_4122);
  not g8028 (n_4123, n4546);
  and g8029 (n4547, n648, n_4123);
  not g8030 (n_4124, n4547);
  and g8031 (n4548, n652, n_4124);
  not g8032 (n_4125, n4548);
  and g8033 (n4549, n656, n_4125);
  not g8034 (n_4126, n4549);
  and g8035 (n4550, n660, n_4126);
  not g8036 (n_4127, n4550);
  and g8037 (n4551, n664, n_4127);
  not g8038 (n_4128, n4551);
  and g8039 (n4552, n668, n_4128);
  not g8040 (n_4129, n4552);
  and g8041 (n4553, n672, n_4129);
  not g8042 (n_4130, n4553);
  and g8043 (n4554, n676, n_4130);
  not g8044 (n_4131, n4554);
  and g8045 (n4555, n680, n_4131);
  not g8046 (n_4132, n4555);
  and g8047 (n4556, n684, n_4132);
  not g8048 (n_4133, n4556);
  and g8049 (n4557, n688, n_4133);
  not g8050 (n_4134, n4557);
  and g8051 (n4558, n692, n_4134);
  not g8052 (n_4135, n4558);
  and g8053 (n4559, n696, n_4135);
  not g8054 (n_4136, n4559);
  and g8055 (n4560, n700, n_4136);
  not g8056 (n_4137, n4560);
  and g8057 (n4561, n704, n_4137);
  not g8058 (n_4138, n4561);
  and g8059 (n4562, n708, n_4138);
  not g8060 (n_4139, n4562);
  and g8061 (n4563, n712, n_4139);
  not g8062 (n_4140, n4563);
  and g8063 (n4564, n716, n_4140);
  not g8064 (n_4141, n4564);
  and g8065 (n4565, n720, n_4141);
  not g8066 (n_4142, n4565);
  and g8067 (n4566, n1484, n_4142);
  not g8068 (n_4143, n4566);
  and g8069 (n4567, n1486, n_4143);
  not g8070 (n_4144, n4567);
  and g8071 (n4568, n1750, n_4144);
  not g8072 (n_4145, n4568);
  and g8073 (n4569, n731, n_4145);
  not g8074 (n_4146, n4569);
  and g8075 (n4570, n735, n_4146);
  not g8076 (n_4147, n4570);
  and g8077 (n4571, n739, n_4147);
  not g8078 (n_4148, n4571);
  and g8079 (n4572, n743, n_4148);
  not g8080 (n_4149, n4572);
  and g8081 (n4573, n747, n_4149);
  not g8082 (n_4150, n4573);
  and g8083 (n4574, n751, n_4150);
  not g8084 (n_4151, n4574);
  and g8085 (n4575, n755, n_4151);
  not g8086 (n_4152, n4575);
  and g8087 (n4576, n759, n_4152);
  not g8088 (n_4153, n4576);
  and g8089 (n4577, n763, n_4153);
  not g8090 (n_4154, n4577);
  and g8091 (n4578, n767, n_4154);
  not g8092 (n_4155, n4578);
  and g8093 (n4579, n771, n_4155);
  not g8094 (n_4156, n4579);
  and g8095 (n4580, n775, n_4156);
  not g8096 (n_4157, n4580);
  and g8097 (n4581, n779, n_4157);
  not g8098 (n_4158, n4581);
  and g8099 (n4582, n783, n_4158);
  not g8100 (n_4159, n4582);
  and g8101 (n4583, n787, n_4159);
  not g8102 (n_4160, n4583);
  and g8103 (n4584, n791, n_4160);
  not g8104 (n_4161, n4584);
  and g8105 (n4585, n795, n_4161);
  not g8106 (n_4162, n4585);
  and g8107 (n4586, n799, n_4162);
  not g8108 (n_4163, n4586);
  and g8109 (n4587, n803, n_4163);
  not g8110 (n_4164, n4587);
  and g8111 (n4588, n807, n_4164);
  not g8112 (n_4165, n4588);
  and g8113 (n4589, n811, n_4165);
  not g8114 (n_4166, n4589);
  and g8115 (n4590, n815, n_4166);
  not g8116 (n_4167, n4590);
  and g8117 (n4591, n819, n_4167);
  and g8118 (n4592, \req[39] , n_671);
  not g8119 (n_4168, n4591);
  and g8120 (\grant[39] , n_4168, n4592);
  not g8121 (n_4169, n1163);
  and g8122 (n4594, n830, n_4169);
  not g8123 (n_4170, n4594);
  and g8124 (n4595, n835, n_4170);
  not g8125 (n_4171, n4595);
  and g8126 (n4596, n839, n_4171);
  not g8127 (n_4172, n4596);
  and g8128 (n4597, n843, n_4172);
  not g8129 (n_4173, n4597);
  and g8130 (n4598, n847, n_4173);
  not g8131 (n_4174, n4598);
  and g8132 (n4599, n851, n_4174);
  not g8133 (n_4175, n4599);
  and g8134 (n4600, n855, n_4175);
  not g8135 (n_4176, n4600);
  and g8136 (n4601, n859, n_4176);
  not g8137 (n_4177, n4601);
  and g8138 (n4602, n863, n_4177);
  not g8139 (n_4178, n4602);
  and g8140 (n4603, n867, n_4178);
  not g8141 (n_4179, n4603);
  and g8142 (n4604, n871, n_4179);
  not g8143 (n_4180, n4604);
  and g8144 (n4605, n875, n_4180);
  not g8145 (n_4181, n4605);
  and g8146 (n4606, n879, n_4181);
  not g8147 (n_4182, n4606);
  and g8148 (n4607, n883, n_4182);
  not g8149 (n_4183, n4607);
  and g8150 (n4608, n887, n_4183);
  not g8151 (n_4184, n4608);
  and g8152 (n4609, n891, n_4184);
  not g8153 (n_4185, n4609);
  and g8154 (n4610, n895, n_4185);
  not g8155 (n_4186, n4610);
  and g8156 (n4611, n899, n_4186);
  not g8157 (n_4187, n4611);
  and g8158 (n4612, n903, n_4187);
  not g8159 (n_4188, n4612);
  and g8160 (n4613, n907, n_4188);
  not g8161 (n_4189, n4613);
  and g8162 (n4614, n911, n_4189);
  not g8163 (n_4190, n4614);
  and g8164 (n4615, n915, n_4190);
  not g8165 (n_4191, n4615);
  and g8166 (n4616, n919, n_4191);
  not g8167 (n_4192, n4616);
  and g8168 (n4617, n923, n_4192);
  not g8169 (n_4193, n4617);
  and g8170 (n4618, n927, n_4193);
  not g8171 (n_4194, n4618);
  and g8172 (n4619, n931, n_4194);
  not g8173 (n_4195, n4619);
  and g8174 (n4620, n935, n_4195);
  not g8175 (n_4196, n4620);
  and g8176 (n4621, n939, n_4196);
  not g8177 (n_4197, n4621);
  and g8178 (n4622, n943, n_4197);
  not g8179 (n_4198, n4622);
  and g8180 (n4623, n947, n_4198);
  not g8181 (n_4199, n4623);
  and g8182 (n4624, n951, n_4199);
  not g8183 (n_4200, n4624);
  and g8184 (n4625, n955, n_4200);
  not g8185 (n_4201, n4625);
  and g8186 (n4626, n959, n_4201);
  not g8187 (n_4202, n4626);
  and g8188 (n4627, n963, n_4202);
  not g8189 (n_4203, n4627);
  and g8190 (n4628, n967, n_4203);
  not g8191 (n_4204, n4628);
  and g8192 (n4629, n971, n_4204);
  not g8193 (n_4205, n4629);
  and g8194 (n4630, n975, n_4205);
  not g8195 (n_4206, n4630);
  and g8196 (n4631, n979, n_4206);
  not g8197 (n_4207, n4631);
  and g8198 (n4632, n983, n_4207);
  not g8199 (n_4208, n4632);
  and g8200 (n4633, n987, n_4208);
  not g8201 (n_4209, n4633);
  and g8202 (n4634, n991, n_4209);
  not g8203 (n_4210, n4634);
  and g8204 (n4635, n995, n_4210);
  not g8205 (n_4211, n4635);
  and g8206 (n4636, n999, n_4211);
  not g8207 (n_4212, n4636);
  and g8208 (n4637, n1003, n_4212);
  not g8209 (n_4213, n4637);
  and g8210 (n4638, n1007, n_4213);
  not g8211 (n_4214, n4638);
  and g8212 (n4639, n1011, n_4214);
  not g8213 (n_4215, n4639);
  and g8214 (n4640, n1015, n_4215);
  not g8215 (n_4216, n4640);
  and g8216 (n4641, n1019, n_4216);
  not g8217 (n_4217, n4641);
  and g8218 (n4642, n1023, n_4217);
  not g8219 (n_4218, n4642);
  and g8220 (n4643, n1027, n_4218);
  not g8221 (n_4219, n4643);
  and g8222 (n4644, n1031, n_4219);
  not g8223 (n_4220, n4644);
  and g8224 (n4645, n1035, n_4220);
  not g8225 (n_4221, n4645);
  and g8226 (n4646, n1039, n_4221);
  not g8227 (n_4222, n4646);
  and g8228 (n4647, n1043, n_4222);
  not g8229 (n_4223, n4647);
  and g8230 (n4648, n1047, n_4223);
  not g8231 (n_4224, n4648);
  and g8232 (n4649, n1051, n_4224);
  not g8233 (n_4225, n4649);
  and g8234 (n4650, n1055, n_4225);
  not g8235 (n_4226, n4650);
  and g8236 (n4651, n1059, n_4226);
  not g8237 (n_4227, n4651);
  and g8238 (n4652, n1574, n_4227);
  not g8239 (n_4228, n4652);
  and g8240 (n4653, n1576, n_4228);
  not g8241 (n_4229, n4653);
  and g8242 (n4654, n1837, n_4229);
  not g8243 (n_4230, n4654);
  and g8244 (n4655, n1068, n_4230);
  not g8245 (n_4231, n4655);
  and g8246 (n4656, n1072, n_4231);
  not g8247 (n_4232, n4656);
  and g8248 (n4657, n1076, n_4232);
  not g8249 (n_4233, n4657);
  and g8250 (n4658, n1080, n_4233);
  not g8251 (n_4234, n4658);
  and g8252 (n4659, n1084, n_4234);
  not g8253 (n_4235, n4659);
  and g8254 (n4660, n1088, n_4235);
  not g8255 (n_4236, n4660);
  and g8256 (n4661, n1092, n_4236);
  not g8257 (n_4237, n4661);
  and g8258 (n4662, n1096, n_4237);
  not g8259 (n_4238, n4662);
  and g8260 (n4663, n1100, n_4238);
  not g8261 (n_4239, n4663);
  and g8262 (n4664, n1104, n_4239);
  not g8263 (n_4240, n4664);
  and g8264 (n4665, n1108, n_4240);
  not g8265 (n_4241, n4665);
  and g8266 (n4666, n1112, n_4241);
  not g8267 (n_4242, n4666);
  and g8268 (n4667, n1116, n_4242);
  not g8269 (n_4243, n4667);
  and g8270 (n4668, n1120, n_4243);
  not g8271 (n_4244, n4668);
  and g8272 (n4669, n1124, n_4244);
  not g8273 (n_4245, n4669);
  and g8274 (n4670, n1128, n_4245);
  not g8275 (n_4246, n4670);
  and g8276 (n4671, n1132, n_4246);
  not g8277 (n_4247, n4671);
  and g8278 (n4672, n1136, n_4247);
  not g8279 (n_4248, n4672);
  and g8280 (n4673, n1140, n_4248);
  not g8281 (n_4249, n4673);
  and g8282 (n4674, n1144, n_4249);
  not g8283 (n_4250, n4674);
  and g8284 (n4675, n1148, n_4250);
  not g8285 (n_4251, n4675);
  and g8286 (n4676, n1152, n_4251);
  not g8287 (n_4252, n4676);
  and g8288 (n4677, n1156, n_4252);
  and g8289 (n4678, \req[40] , n_899);
  not g8290 (n_4253, n4677);
  and g8291 (\grant[40] , n_4253, n4678);
  not g8292 (n_4254, n495);
  and g8293 (n4680, n_4254, n1167);
  not g8294 (n_4255, n4680);
  and g8295 (n4681, n1172, n_4255);
  not g8296 (n_4256, n4681);
  and g8297 (n4682, n1176, n_4256);
  not g8298 (n_4257, n4682);
  and g8299 (n4683, n1180, n_4257);
  not g8300 (n_4258, n4683);
  and g8301 (n4684, n1184, n_4258);
  not g8302 (n_4259, n4684);
  and g8303 (n4685, n1188, n_4259);
  not g8304 (n_4260, n4685);
  and g8305 (n4686, n1192, n_4260);
  not g8306 (n_4261, n4686);
  and g8307 (n4687, n1196, n_4261);
  not g8308 (n_4262, n4687);
  and g8309 (n4688, n1200, n_4262);
  not g8310 (n_4263, n4688);
  and g8311 (n4689, n1204, n_4263);
  not g8312 (n_4264, n4689);
  and g8313 (n4690, n1208, n_4264);
  not g8314 (n_4265, n4690);
  and g8315 (n4691, n1212, n_4265);
  not g8316 (n_4266, n4691);
  and g8317 (n4692, n1216, n_4266);
  not g8318 (n_4267, n4692);
  and g8319 (n4693, n1220, n_4267);
  not g8320 (n_4268, n4693);
  and g8321 (n4694, n1224, n_4268);
  not g8322 (n_4269, n4694);
  and g8323 (n4695, n1228, n_4269);
  not g8324 (n_4270, n4695);
  and g8325 (n4696, n1232, n_4270);
  not g8326 (n_4271, n4696);
  and g8327 (n4697, n1236, n_4271);
  not g8328 (n_4272, n4697);
  and g8329 (n4698, n1240, n_4272);
  not g8330 (n_4273, n4698);
  and g8331 (n4699, n1244, n_4273);
  not g8332 (n_4274, n4699);
  and g8333 (n4700, n1248, n_4274);
  not g8334 (n_4275, n4700);
  and g8335 (n4701, n1252, n_4275);
  not g8336 (n_4276, n4701);
  and g8337 (n4702, n1256, n_4276);
  not g8338 (n_4277, n4702);
  and g8339 (n4703, n1260, n_4277);
  not g8340 (n_4278, n4703);
  and g8341 (n4704, n1264, n_4278);
  not g8342 (n_4279, n4704);
  and g8343 (n4705, n1268, n_4279);
  not g8344 (n_4280, n4705);
  and g8345 (n4706, n1272, n_4280);
  not g8346 (n_4281, n4706);
  and g8347 (n4707, n1276, n_4281);
  not g8348 (n_4282, n4707);
  and g8349 (n4708, n1280, n_4282);
  not g8350 (n_4283, n4708);
  and g8351 (n4709, n1284, n_4283);
  not g8352 (n_4284, n4709);
  and g8353 (n4710, n1288, n_4284);
  not g8354 (n_4285, n4710);
  and g8355 (n4711, n1292, n_4285);
  not g8356 (n_4286, n4711);
  and g8357 (n4712, n1296, n_4286);
  not g8358 (n_4287, n4712);
  and g8359 (n4713, n1300, n_4287);
  not g8360 (n_4288, n4713);
  and g8361 (n4714, n1304, n_4288);
  not g8362 (n_4289, n4714);
  and g8363 (n4715, n1308, n_4289);
  not g8364 (n_4290, n4715);
  and g8365 (n4716, n1312, n_4290);
  not g8366 (n_4291, n4716);
  and g8367 (n4717, n1316, n_4291);
  not g8368 (n_4292, n4717);
  and g8369 (n4718, n1320, n_4292);
  not g8370 (n_4293, n4718);
  and g8371 (n4719, n1324, n_4293);
  not g8372 (n_4294, n4719);
  and g8373 (n4720, n1328, n_4294);
  not g8374 (n_4295, n4720);
  and g8375 (n4721, n1332, n_4295);
  not g8376 (n_4296, n4721);
  and g8377 (n4722, n1336, n_4296);
  not g8378 (n_4297, n4722);
  and g8379 (n4723, n1340, n_4297);
  not g8380 (n_4298, n4723);
  and g8381 (n4724, n1344, n_4298);
  not g8382 (n_4299, n4724);
  and g8383 (n4725, n1348, n_4299);
  not g8384 (n_4300, n4725);
  and g8385 (n4726, n1352, n_4300);
  not g8386 (n_4301, n4726);
  and g8387 (n4727, n1356, n_4301);
  not g8388 (n_4302, n4727);
  and g8389 (n4728, n1360, n_4302);
  not g8390 (n_4303, n4728);
  and g8391 (n4729, n1364, n_4303);
  not g8392 (n_4304, n4729);
  and g8393 (n4730, n1368, n_4304);
  not g8394 (n_4305, n4730);
  and g8395 (n4731, n1372, n_4305);
  not g8396 (n_4306, n4731);
  and g8397 (n4732, n1376, n_4306);
  not g8398 (n_4307, n4732);
  and g8399 (n4733, n1380, n_4307);
  not g8400 (n_4308, n4733);
  and g8401 (n4734, n1384, n_4308);
  not g8402 (n_4309, n4734);
  and g8403 (n4735, n1388, n_4309);
  not g8404 (n_4310, n4735);
  and g8405 (n4736, n1392, n_4310);
  not g8406 (n_4311, n4736);
  and g8407 (n4737, n1396, n_4311);
  not g8408 (n_4312, n4737);
  and g8409 (n4738, n1663, n_4312);
  not g8410 (n_4313, n4738);
  and g8411 (n4739, n392, n_4313);
  not g8412 (n_4314, n4739);
  and g8413 (n4740, n396, n_4314);
  not g8414 (n_4315, n4740);
  and g8415 (n4741, n400, n_4315);
  not g8416 (n_4316, n4741);
  and g8417 (n4742, n404, n_4316);
  not g8418 (n_4317, n4742);
  and g8419 (n4743, n408, n_4317);
  not g8420 (n_4318, n4743);
  and g8421 (n4744, n412, n_4318);
  not g8422 (n_4319, n4744);
  and g8423 (n4745, n416, n_4319);
  not g8424 (n_4320, n4745);
  and g8425 (n4746, n420, n_4320);
  not g8426 (n_4321, n4746);
  and g8427 (n4747, n424, n_4321);
  not g8428 (n_4322, n4747);
  and g8429 (n4748, n428, n_4322);
  not g8430 (n_4323, n4748);
  and g8431 (n4749, n432, n_4323);
  not g8432 (n_4324, n4749);
  and g8433 (n4750, n436, n_4324);
  not g8434 (n_4325, n4750);
  and g8435 (n4751, n440, n_4325);
  not g8436 (n_4326, n4751);
  and g8437 (n4752, n444, n_4326);
  not g8438 (n_4327, n4752);
  and g8439 (n4753, n448, n_4327);
  not g8440 (n_4328, n4753);
  and g8441 (n4754, n452, n_4328);
  not g8442 (n_4329, n4754);
  and g8443 (n4755, n456, n_4329);
  not g8444 (n_4330, n4755);
  and g8445 (n4756, n460, n_4330);
  not g8446 (n_4331, n4756);
  and g8447 (n4757, n464, n_4331);
  not g8448 (n_4332, n4757);
  and g8449 (n4758, n468, n_4332);
  not g8450 (n_4333, n4758);
  and g8451 (n4759, n472, n_4333);
  not g8452 (n_4334, n4759);
  and g8453 (n4760, n476, n_4334);
  not g8454 (n_4335, n4760);
  and g8455 (n4761, n480, n_4335);
  not g8456 (n_4336, n4761);
  and g8457 (n4762, n484, n_4336);
  not g8458 (n_4337, n4762);
  and g8459 (n4763, n488, n_4337);
  and g8460 (n4764, \req[41] , n_192);
  not g8461 (n_4338, n4763);
  and g8462 (\grant[41] , n_4338, n4764);
  not g8463 (n_4339, n834);
  and g8464 (n4766, n499, n_4339);
  not g8465 (n_4340, n4766);
  and g8466 (n4767, n504, n_4340);
  not g8467 (n_4341, n4767);
  and g8468 (n4768, n508, n_4341);
  not g8469 (n_4342, n4768);
  and g8470 (n4769, n512, n_4342);
  not g8471 (n_4343, n4769);
  and g8472 (n4770, n516, n_4343);
  not g8473 (n_4344, n4770);
  and g8474 (n4771, n520, n_4344);
  not g8475 (n_4345, n4771);
  and g8476 (n4772, n524, n_4345);
  not g8477 (n_4346, n4772);
  and g8478 (n4773, n528, n_4346);
  not g8479 (n_4347, n4773);
  and g8480 (n4774, n532, n_4347);
  not g8481 (n_4348, n4774);
  and g8482 (n4775, n536, n_4348);
  not g8483 (n_4349, n4775);
  and g8484 (n4776, n540, n_4349);
  not g8485 (n_4350, n4776);
  and g8486 (n4777, n544, n_4350);
  not g8487 (n_4351, n4777);
  and g8488 (n4778, n548, n_4351);
  not g8489 (n_4352, n4778);
  and g8490 (n4779, n552, n_4352);
  not g8491 (n_4353, n4779);
  and g8492 (n4780, n556, n_4353);
  not g8493 (n_4354, n4780);
  and g8494 (n4781, n560, n_4354);
  not g8495 (n_4355, n4781);
  and g8496 (n4782, n564, n_4355);
  not g8497 (n_4356, n4782);
  and g8498 (n4783, n568, n_4356);
  not g8499 (n_4357, n4783);
  and g8500 (n4784, n572, n_4357);
  not g8501 (n_4358, n4784);
  and g8502 (n4785, n576, n_4358);
  not g8503 (n_4359, n4785);
  and g8504 (n4786, n580, n_4359);
  not g8505 (n_4360, n4786);
  and g8506 (n4787, n584, n_4360);
  not g8507 (n_4361, n4787);
  and g8508 (n4788, n588, n_4361);
  not g8509 (n_4362, n4788);
  and g8510 (n4789, n592, n_4362);
  not g8511 (n_4363, n4789);
  and g8512 (n4790, n596, n_4363);
  not g8513 (n_4364, n4790);
  and g8514 (n4791, n600, n_4364);
  not g8515 (n_4365, n4791);
  and g8516 (n4792, n604, n_4365);
  not g8517 (n_4366, n4792);
  and g8518 (n4793, n608, n_4366);
  not g8519 (n_4367, n4793);
  and g8520 (n4794, n612, n_4367);
  not g8521 (n_4368, n4794);
  and g8522 (n4795, n616, n_4368);
  not g8523 (n_4369, n4795);
  and g8524 (n4796, n620, n_4369);
  not g8525 (n_4370, n4796);
  and g8526 (n4797, n624, n_4370);
  not g8527 (n_4371, n4797);
  and g8528 (n4798, n628, n_4371);
  not g8529 (n_4372, n4798);
  and g8530 (n4799, n632, n_4372);
  not g8531 (n_4373, n4799);
  and g8532 (n4800, n636, n_4373);
  not g8533 (n_4374, n4800);
  and g8534 (n4801, n640, n_4374);
  not g8535 (n_4375, n4801);
  and g8536 (n4802, n644, n_4375);
  not g8537 (n_4376, n4802);
  and g8538 (n4803, n648, n_4376);
  not g8539 (n_4377, n4803);
  and g8540 (n4804, n652, n_4377);
  not g8541 (n_4378, n4804);
  and g8542 (n4805, n656, n_4378);
  not g8543 (n_4379, n4805);
  and g8544 (n4806, n660, n_4379);
  not g8545 (n_4380, n4806);
  and g8546 (n4807, n664, n_4380);
  not g8547 (n_4381, n4807);
  and g8548 (n4808, n668, n_4381);
  not g8549 (n_4382, n4808);
  and g8550 (n4809, n672, n_4382);
  not g8551 (n_4383, n4809);
  and g8552 (n4810, n676, n_4383);
  not g8553 (n_4384, n4810);
  and g8554 (n4811, n680, n_4384);
  not g8555 (n_4385, n4811);
  and g8556 (n4812, n684, n_4385);
  not g8557 (n_4386, n4812);
  and g8558 (n4813, n688, n_4386);
  not g8559 (n_4387, n4813);
  and g8560 (n4814, n692, n_4387);
  not g8561 (n_4388, n4814);
  and g8562 (n4815, n696, n_4388);
  not g8563 (n_4389, n4815);
  and g8564 (n4816, n700, n_4389);
  not g8565 (n_4390, n4816);
  and g8566 (n4817, n704, n_4390);
  not g8567 (n_4391, n4817);
  and g8568 (n4818, n708, n_4391);
  not g8569 (n_4392, n4818);
  and g8570 (n4819, n712, n_4392);
  not g8571 (n_4393, n4819);
  and g8572 (n4820, n716, n_4393);
  not g8573 (n_4394, n4820);
  and g8574 (n4821, n720, n_4394);
  not g8575 (n_4395, n4821);
  and g8576 (n4822, n1484, n_4395);
  not g8577 (n_4396, n4822);
  and g8578 (n4823, n1486, n_4396);
  not g8579 (n_4397, n4823);
  and g8580 (n4824, n1750, n_4397);
  not g8581 (n_4398, n4824);
  and g8582 (n4825, n731, n_4398);
  not g8583 (n_4399, n4825);
  and g8584 (n4826, n735, n_4399);
  not g8585 (n_4400, n4826);
  and g8586 (n4827, n739, n_4400);
  not g8587 (n_4401, n4827);
  and g8588 (n4828, n743, n_4401);
  not g8589 (n_4402, n4828);
  and g8590 (n4829, n747, n_4402);
  not g8591 (n_4403, n4829);
  and g8592 (n4830, n751, n_4403);
  not g8593 (n_4404, n4830);
  and g8594 (n4831, n755, n_4404);
  not g8595 (n_4405, n4831);
  and g8596 (n4832, n759, n_4405);
  not g8597 (n_4406, n4832);
  and g8598 (n4833, n763, n_4406);
  not g8599 (n_4407, n4833);
  and g8600 (n4834, n767, n_4407);
  not g8601 (n_4408, n4834);
  and g8602 (n4835, n771, n_4408);
  not g8603 (n_4409, n4835);
  and g8604 (n4836, n775, n_4409);
  not g8605 (n_4410, n4836);
  and g8606 (n4837, n779, n_4410);
  not g8607 (n_4411, n4837);
  and g8608 (n4838, n783, n_4411);
  not g8609 (n_4412, n4838);
  and g8610 (n4839, n787, n_4412);
  not g8611 (n_4413, n4839);
  and g8612 (n4840, n791, n_4413);
  not g8613 (n_4414, n4840);
  and g8614 (n4841, n795, n_4414);
  not g8615 (n_4415, n4841);
  and g8616 (n4842, n799, n_4415);
  not g8617 (n_4416, n4842);
  and g8618 (n4843, n803, n_4416);
  not g8619 (n_4417, n4843);
  and g8620 (n4844, n807, n_4417);
  not g8621 (n_4418, n4844);
  and g8622 (n4845, n811, n_4418);
  not g8623 (n_4419, n4845);
  and g8624 (n4846, n815, n_4419);
  not g8625 (n_4420, n4846);
  and g8626 (n4847, n819, n_4420);
  not g8627 (n_4421, n4847);
  and g8628 (n4848, n823, n_4421);
  not g8629 (n_4422, n4848);
  and g8630 (n4849, n827, n_4422);
  and g8631 (n4850, \req[42] , n_677);
  not g8632 (n_4423, n4849);
  and g8633 (\grant[42] , n_4423, n4850);
  not g8634 (n_4424, n1171);
  and g8635 (n4852, n838, n_4424);
  not g8636 (n_4425, n4852);
  and g8637 (n4853, n843, n_4425);
  not g8638 (n_4426, n4853);
  and g8639 (n4854, n847, n_4426);
  not g8640 (n_4427, n4854);
  and g8641 (n4855, n851, n_4427);
  not g8642 (n_4428, n4855);
  and g8643 (n4856, n855, n_4428);
  not g8644 (n_4429, n4856);
  and g8645 (n4857, n859, n_4429);
  not g8646 (n_4430, n4857);
  and g8647 (n4858, n863, n_4430);
  not g8648 (n_4431, n4858);
  and g8649 (n4859, n867, n_4431);
  not g8650 (n_4432, n4859);
  and g8651 (n4860, n871, n_4432);
  not g8652 (n_4433, n4860);
  and g8653 (n4861, n875, n_4433);
  not g8654 (n_4434, n4861);
  and g8655 (n4862, n879, n_4434);
  not g8656 (n_4435, n4862);
  and g8657 (n4863, n883, n_4435);
  not g8658 (n_4436, n4863);
  and g8659 (n4864, n887, n_4436);
  not g8660 (n_4437, n4864);
  and g8661 (n4865, n891, n_4437);
  not g8662 (n_4438, n4865);
  and g8663 (n4866, n895, n_4438);
  not g8664 (n_4439, n4866);
  and g8665 (n4867, n899, n_4439);
  not g8666 (n_4440, n4867);
  and g8667 (n4868, n903, n_4440);
  not g8668 (n_4441, n4868);
  and g8669 (n4869, n907, n_4441);
  not g8670 (n_4442, n4869);
  and g8671 (n4870, n911, n_4442);
  not g8672 (n_4443, n4870);
  and g8673 (n4871, n915, n_4443);
  not g8674 (n_4444, n4871);
  and g8675 (n4872, n919, n_4444);
  not g8676 (n_4445, n4872);
  and g8677 (n4873, n923, n_4445);
  not g8678 (n_4446, n4873);
  and g8679 (n4874, n927, n_4446);
  not g8680 (n_4447, n4874);
  and g8681 (n4875, n931, n_4447);
  not g8682 (n_4448, n4875);
  and g8683 (n4876, n935, n_4448);
  not g8684 (n_4449, n4876);
  and g8685 (n4877, n939, n_4449);
  not g8686 (n_4450, n4877);
  and g8687 (n4878, n943, n_4450);
  not g8688 (n_4451, n4878);
  and g8689 (n4879, n947, n_4451);
  not g8690 (n_4452, n4879);
  and g8691 (n4880, n951, n_4452);
  not g8692 (n_4453, n4880);
  and g8693 (n4881, n955, n_4453);
  not g8694 (n_4454, n4881);
  and g8695 (n4882, n959, n_4454);
  not g8696 (n_4455, n4882);
  and g8697 (n4883, n963, n_4455);
  not g8698 (n_4456, n4883);
  and g8699 (n4884, n967, n_4456);
  not g8700 (n_4457, n4884);
  and g8701 (n4885, n971, n_4457);
  not g8702 (n_4458, n4885);
  and g8703 (n4886, n975, n_4458);
  not g8704 (n_4459, n4886);
  and g8705 (n4887, n979, n_4459);
  not g8706 (n_4460, n4887);
  and g8707 (n4888, n983, n_4460);
  not g8708 (n_4461, n4888);
  and g8709 (n4889, n987, n_4461);
  not g8710 (n_4462, n4889);
  and g8711 (n4890, n991, n_4462);
  not g8712 (n_4463, n4890);
  and g8713 (n4891, n995, n_4463);
  not g8714 (n_4464, n4891);
  and g8715 (n4892, n999, n_4464);
  not g8716 (n_4465, n4892);
  and g8717 (n4893, n1003, n_4465);
  not g8718 (n_4466, n4893);
  and g8719 (n4894, n1007, n_4466);
  not g8720 (n_4467, n4894);
  and g8721 (n4895, n1011, n_4467);
  not g8722 (n_4468, n4895);
  and g8723 (n4896, n1015, n_4468);
  not g8724 (n_4469, n4896);
  and g8725 (n4897, n1019, n_4469);
  not g8726 (n_4470, n4897);
  and g8727 (n4898, n1023, n_4470);
  not g8728 (n_4471, n4898);
  and g8729 (n4899, n1027, n_4471);
  not g8730 (n_4472, n4899);
  and g8731 (n4900, n1031, n_4472);
  not g8732 (n_4473, n4900);
  and g8733 (n4901, n1035, n_4473);
  not g8734 (n_4474, n4901);
  and g8735 (n4902, n1039, n_4474);
  not g8736 (n_4475, n4902);
  and g8737 (n4903, n1043, n_4475);
  not g8738 (n_4476, n4903);
  and g8739 (n4904, n1047, n_4476);
  not g8740 (n_4477, n4904);
  and g8741 (n4905, n1051, n_4477);
  not g8742 (n_4478, n4905);
  and g8743 (n4906, n1055, n_4478);
  not g8744 (n_4479, n4906);
  and g8745 (n4907, n1059, n_4479);
  not g8746 (n_4480, n4907);
  and g8747 (n4908, n1574, n_4480);
  not g8748 (n_4481, n4908);
  and g8749 (n4909, n1576, n_4481);
  not g8750 (n_4482, n4909);
  and g8751 (n4910, n1837, n_4482);
  not g8752 (n_4483, n4910);
  and g8753 (n4911, n1068, n_4483);
  not g8754 (n_4484, n4911);
  and g8755 (n4912, n1072, n_4484);
  not g8756 (n_4485, n4912);
  and g8757 (n4913, n1076, n_4485);
  not g8758 (n_4486, n4913);
  and g8759 (n4914, n1080, n_4486);
  not g8760 (n_4487, n4914);
  and g8761 (n4915, n1084, n_4487);
  not g8762 (n_4488, n4915);
  and g8763 (n4916, n1088, n_4488);
  not g8764 (n_4489, n4916);
  and g8765 (n4917, n1092, n_4489);
  not g8766 (n_4490, n4917);
  and g8767 (n4918, n1096, n_4490);
  not g8768 (n_4491, n4918);
  and g8769 (n4919, n1100, n_4491);
  not g8770 (n_4492, n4919);
  and g8771 (n4920, n1104, n_4492);
  not g8772 (n_4493, n4920);
  and g8773 (n4921, n1108, n_4493);
  not g8774 (n_4494, n4921);
  and g8775 (n4922, n1112, n_4494);
  not g8776 (n_4495, n4922);
  and g8777 (n4923, n1116, n_4495);
  not g8778 (n_4496, n4923);
  and g8779 (n4924, n1120, n_4496);
  not g8780 (n_4497, n4924);
  and g8781 (n4925, n1124, n_4497);
  not g8782 (n_4498, n4925);
  and g8783 (n4926, n1128, n_4498);
  not g8784 (n_4499, n4926);
  and g8785 (n4927, n1132, n_4499);
  not g8786 (n_4500, n4927);
  and g8787 (n4928, n1136, n_4500);
  not g8788 (n_4501, n4928);
  and g8789 (n4929, n1140, n_4501);
  not g8790 (n_4502, n4929);
  and g8791 (n4930, n1144, n_4502);
  not g8792 (n_4503, n4930);
  and g8793 (n4931, n1148, n_4503);
  not g8794 (n_4504, n4931);
  and g8795 (n4932, n1152, n_4504);
  not g8796 (n_4505, n4932);
  and g8797 (n4933, n1156, n_4505);
  not g8798 (n_4506, n4933);
  and g8799 (n4934, n1160, n_4506);
  not g8800 (n_4507, n4934);
  and g8801 (n4935, n1164, n_4507);
  and g8802 (n4936, \req[43] , n_903);
  not g8803 (n_4508, n4935);
  and g8804 (\grant[43] , n_4508, n4936);
  not g8805 (n_4509, n503);
  and g8806 (n4938, n_4509, n1175);
  not g8807 (n_4510, n4938);
  and g8808 (n4939, n1180, n_4510);
  not g8809 (n_4511, n4939);
  and g8810 (n4940, n1184, n_4511);
  not g8811 (n_4512, n4940);
  and g8812 (n4941, n1188, n_4512);
  not g8813 (n_4513, n4941);
  and g8814 (n4942, n1192, n_4513);
  not g8815 (n_4514, n4942);
  and g8816 (n4943, n1196, n_4514);
  not g8817 (n_4515, n4943);
  and g8818 (n4944, n1200, n_4515);
  not g8819 (n_4516, n4944);
  and g8820 (n4945, n1204, n_4516);
  not g8821 (n_4517, n4945);
  and g8822 (n4946, n1208, n_4517);
  not g8823 (n_4518, n4946);
  and g8824 (n4947, n1212, n_4518);
  not g8825 (n_4519, n4947);
  and g8826 (n4948, n1216, n_4519);
  not g8827 (n_4520, n4948);
  and g8828 (n4949, n1220, n_4520);
  not g8829 (n_4521, n4949);
  and g8830 (n4950, n1224, n_4521);
  not g8831 (n_4522, n4950);
  and g8832 (n4951, n1228, n_4522);
  not g8833 (n_4523, n4951);
  and g8834 (n4952, n1232, n_4523);
  not g8835 (n_4524, n4952);
  and g8836 (n4953, n1236, n_4524);
  not g8837 (n_4525, n4953);
  and g8838 (n4954, n1240, n_4525);
  not g8839 (n_4526, n4954);
  and g8840 (n4955, n1244, n_4526);
  not g8841 (n_4527, n4955);
  and g8842 (n4956, n1248, n_4527);
  not g8843 (n_4528, n4956);
  and g8844 (n4957, n1252, n_4528);
  not g8845 (n_4529, n4957);
  and g8846 (n4958, n1256, n_4529);
  not g8847 (n_4530, n4958);
  and g8848 (n4959, n1260, n_4530);
  not g8849 (n_4531, n4959);
  and g8850 (n4960, n1264, n_4531);
  not g8851 (n_4532, n4960);
  and g8852 (n4961, n1268, n_4532);
  not g8853 (n_4533, n4961);
  and g8854 (n4962, n1272, n_4533);
  not g8855 (n_4534, n4962);
  and g8856 (n4963, n1276, n_4534);
  not g8857 (n_4535, n4963);
  and g8858 (n4964, n1280, n_4535);
  not g8859 (n_4536, n4964);
  and g8860 (n4965, n1284, n_4536);
  not g8861 (n_4537, n4965);
  and g8862 (n4966, n1288, n_4537);
  not g8863 (n_4538, n4966);
  and g8864 (n4967, n1292, n_4538);
  not g8865 (n_4539, n4967);
  and g8866 (n4968, n1296, n_4539);
  not g8867 (n_4540, n4968);
  and g8868 (n4969, n1300, n_4540);
  not g8869 (n_4541, n4969);
  and g8870 (n4970, n1304, n_4541);
  not g8871 (n_4542, n4970);
  and g8872 (n4971, n1308, n_4542);
  not g8873 (n_4543, n4971);
  and g8874 (n4972, n1312, n_4543);
  not g8875 (n_4544, n4972);
  and g8876 (n4973, n1316, n_4544);
  not g8877 (n_4545, n4973);
  and g8878 (n4974, n1320, n_4545);
  not g8879 (n_4546, n4974);
  and g8880 (n4975, n1324, n_4546);
  not g8881 (n_4547, n4975);
  and g8882 (n4976, n1328, n_4547);
  not g8883 (n_4548, n4976);
  and g8884 (n4977, n1332, n_4548);
  not g8885 (n_4549, n4977);
  and g8886 (n4978, n1336, n_4549);
  not g8887 (n_4550, n4978);
  and g8888 (n4979, n1340, n_4550);
  not g8889 (n_4551, n4979);
  and g8890 (n4980, n1344, n_4551);
  not g8891 (n_4552, n4980);
  and g8892 (n4981, n1348, n_4552);
  not g8893 (n_4553, n4981);
  and g8894 (n4982, n1352, n_4553);
  not g8895 (n_4554, n4982);
  and g8896 (n4983, n1356, n_4554);
  not g8897 (n_4555, n4983);
  and g8898 (n4984, n1360, n_4555);
  not g8899 (n_4556, n4984);
  and g8900 (n4985, n1364, n_4556);
  not g8901 (n_4557, n4985);
  and g8902 (n4986, n1368, n_4557);
  not g8903 (n_4558, n4986);
  and g8904 (n4987, n1372, n_4558);
  not g8905 (n_4559, n4987);
  and g8906 (n4988, n1376, n_4559);
  not g8907 (n_4560, n4988);
  and g8908 (n4989, n1380, n_4560);
  not g8909 (n_4561, n4989);
  and g8910 (n4990, n1384, n_4561);
  not g8911 (n_4562, n4990);
  and g8912 (n4991, n1388, n_4562);
  not g8913 (n_4563, n4991);
  and g8914 (n4992, n1392, n_4563);
  not g8915 (n_4564, n4992);
  and g8916 (n4993, n1396, n_4564);
  not g8917 (n_4565, n4993);
  and g8918 (n4994, n1663, n_4565);
  not g8919 (n_4566, n4994);
  and g8920 (n4995, n392, n_4566);
  not g8921 (n_4567, n4995);
  and g8922 (n4996, n396, n_4567);
  not g8923 (n_4568, n4996);
  and g8924 (n4997, n400, n_4568);
  not g8925 (n_4569, n4997);
  and g8926 (n4998, n404, n_4569);
  not g8927 (n_4570, n4998);
  and g8928 (n4999, n408, n_4570);
  not g8929 (n_4571, n4999);
  and g8930 (n5000, n412, n_4571);
  not g8931 (n_4572, n5000);
  and g8932 (n5001, n416, n_4572);
  not g8933 (n_4573, n5001);
  and g8934 (n5002, n420, n_4573);
  not g8935 (n_4574, n5002);
  and g8936 (n5003, n424, n_4574);
  not g8937 (n_4575, n5003);
  and g8938 (n5004, n428, n_4575);
  not g8939 (n_4576, n5004);
  and g8940 (n5005, n432, n_4576);
  not g8941 (n_4577, n5005);
  and g8942 (n5006, n436, n_4577);
  not g8943 (n_4578, n5006);
  and g8944 (n5007, n440, n_4578);
  not g8945 (n_4579, n5007);
  and g8946 (n5008, n444, n_4579);
  not g8947 (n_4580, n5008);
  and g8948 (n5009, n448, n_4580);
  not g8949 (n_4581, n5009);
  and g8950 (n5010, n452, n_4581);
  not g8951 (n_4582, n5010);
  and g8952 (n5011, n456, n_4582);
  not g8953 (n_4583, n5011);
  and g8954 (n5012, n460, n_4583);
  not g8955 (n_4584, n5012);
  and g8956 (n5013, n464, n_4584);
  not g8957 (n_4585, n5013);
  and g8958 (n5014, n468, n_4585);
  not g8959 (n_4586, n5014);
  and g8960 (n5015, n472, n_4586);
  not g8961 (n_4587, n5015);
  and g8962 (n5016, n476, n_4587);
  not g8963 (n_4588, n5016);
  and g8964 (n5017, n480, n_4588);
  not g8965 (n_4589, n5017);
  and g8966 (n5018, n484, n_4589);
  not g8967 (n_4590, n5018);
  and g8968 (n5019, n488, n_4590);
  not g8969 (n_4591, n5019);
  and g8970 (n5020, n492, n_4591);
  not g8971 (n_4592, n5020);
  and g8972 (n5021, n496, n_4592);
  and g8973 (n5022, \req[44] , n_206);
  not g8974 (n_4593, n5021);
  and g8975 (\grant[44] , n_4593, n5022);
  not g8976 (n_4594, n842);
  and g8977 (n5024, n507, n_4594);
  not g8978 (n_4595, n5024);
  and g8979 (n5025, n512, n_4595);
  not g8980 (n_4596, n5025);
  and g8981 (n5026, n516, n_4596);
  not g8982 (n_4597, n5026);
  and g8983 (n5027, n520, n_4597);
  not g8984 (n_4598, n5027);
  and g8985 (n5028, n524, n_4598);
  not g8986 (n_4599, n5028);
  and g8987 (n5029, n528, n_4599);
  not g8988 (n_4600, n5029);
  and g8989 (n5030, n532, n_4600);
  not g8990 (n_4601, n5030);
  and g8991 (n5031, n536, n_4601);
  not g8992 (n_4602, n5031);
  and g8993 (n5032, n540, n_4602);
  not g8994 (n_4603, n5032);
  and g8995 (n5033, n544, n_4603);
  not g8996 (n_4604, n5033);
  and g8997 (n5034, n548, n_4604);
  not g8998 (n_4605, n5034);
  and g8999 (n5035, n552, n_4605);
  not g9000 (n_4606, n5035);
  and g9001 (n5036, n556, n_4606);
  not g9002 (n_4607, n5036);
  and g9003 (n5037, n560, n_4607);
  not g9004 (n_4608, n5037);
  and g9005 (n5038, n564, n_4608);
  not g9006 (n_4609, n5038);
  and g9007 (n5039, n568, n_4609);
  not g9008 (n_4610, n5039);
  and g9009 (n5040, n572, n_4610);
  not g9010 (n_4611, n5040);
  and g9011 (n5041, n576, n_4611);
  not g9012 (n_4612, n5041);
  and g9013 (n5042, n580, n_4612);
  not g9014 (n_4613, n5042);
  and g9015 (n5043, n584, n_4613);
  not g9016 (n_4614, n5043);
  and g9017 (n5044, n588, n_4614);
  not g9018 (n_4615, n5044);
  and g9019 (n5045, n592, n_4615);
  not g9020 (n_4616, n5045);
  and g9021 (n5046, n596, n_4616);
  not g9022 (n_4617, n5046);
  and g9023 (n5047, n600, n_4617);
  not g9024 (n_4618, n5047);
  and g9025 (n5048, n604, n_4618);
  not g9026 (n_4619, n5048);
  and g9027 (n5049, n608, n_4619);
  not g9028 (n_4620, n5049);
  and g9029 (n5050, n612, n_4620);
  not g9030 (n_4621, n5050);
  and g9031 (n5051, n616, n_4621);
  not g9032 (n_4622, n5051);
  and g9033 (n5052, n620, n_4622);
  not g9034 (n_4623, n5052);
  and g9035 (n5053, n624, n_4623);
  not g9036 (n_4624, n5053);
  and g9037 (n5054, n628, n_4624);
  not g9038 (n_4625, n5054);
  and g9039 (n5055, n632, n_4625);
  not g9040 (n_4626, n5055);
  and g9041 (n5056, n636, n_4626);
  not g9042 (n_4627, n5056);
  and g9043 (n5057, n640, n_4627);
  not g9044 (n_4628, n5057);
  and g9045 (n5058, n644, n_4628);
  not g9046 (n_4629, n5058);
  and g9047 (n5059, n648, n_4629);
  not g9048 (n_4630, n5059);
  and g9049 (n5060, n652, n_4630);
  not g9050 (n_4631, n5060);
  and g9051 (n5061, n656, n_4631);
  not g9052 (n_4632, n5061);
  and g9053 (n5062, n660, n_4632);
  not g9054 (n_4633, n5062);
  and g9055 (n5063, n664, n_4633);
  not g9056 (n_4634, n5063);
  and g9057 (n5064, n668, n_4634);
  not g9058 (n_4635, n5064);
  and g9059 (n5065, n672, n_4635);
  not g9060 (n_4636, n5065);
  and g9061 (n5066, n676, n_4636);
  not g9062 (n_4637, n5066);
  and g9063 (n5067, n680, n_4637);
  not g9064 (n_4638, n5067);
  and g9065 (n5068, n684, n_4638);
  not g9066 (n_4639, n5068);
  and g9067 (n5069, n688, n_4639);
  not g9068 (n_4640, n5069);
  and g9069 (n5070, n692, n_4640);
  not g9070 (n_4641, n5070);
  and g9071 (n5071, n696, n_4641);
  not g9072 (n_4642, n5071);
  and g9073 (n5072, n700, n_4642);
  not g9074 (n_4643, n5072);
  and g9075 (n5073, n704, n_4643);
  not g9076 (n_4644, n5073);
  and g9077 (n5074, n708, n_4644);
  not g9078 (n_4645, n5074);
  and g9079 (n5075, n712, n_4645);
  not g9080 (n_4646, n5075);
  and g9081 (n5076, n716, n_4646);
  not g9082 (n_4647, n5076);
  and g9083 (n5077, n720, n_4647);
  not g9084 (n_4648, n5077);
  and g9085 (n5078, n1484, n_4648);
  not g9086 (n_4649, n5078);
  and g9087 (n5079, n1486, n_4649);
  not g9088 (n_4650, n5079);
  and g9089 (n5080, n1750, n_4650);
  not g9090 (n_4651, n5080);
  and g9091 (n5081, n731, n_4651);
  not g9092 (n_4652, n5081);
  and g9093 (n5082, n735, n_4652);
  not g9094 (n_4653, n5082);
  and g9095 (n5083, n739, n_4653);
  not g9096 (n_4654, n5083);
  and g9097 (n5084, n743, n_4654);
  not g9098 (n_4655, n5084);
  and g9099 (n5085, n747, n_4655);
  not g9100 (n_4656, n5085);
  and g9101 (n5086, n751, n_4656);
  not g9102 (n_4657, n5086);
  and g9103 (n5087, n755, n_4657);
  not g9104 (n_4658, n5087);
  and g9105 (n5088, n759, n_4658);
  not g9106 (n_4659, n5088);
  and g9107 (n5089, n763, n_4659);
  not g9108 (n_4660, n5089);
  and g9109 (n5090, n767, n_4660);
  not g9110 (n_4661, n5090);
  and g9111 (n5091, n771, n_4661);
  not g9112 (n_4662, n5091);
  and g9113 (n5092, n775, n_4662);
  not g9114 (n_4663, n5092);
  and g9115 (n5093, n779, n_4663);
  not g9116 (n_4664, n5093);
  and g9117 (n5094, n783, n_4664);
  not g9118 (n_4665, n5094);
  and g9119 (n5095, n787, n_4665);
  not g9120 (n_4666, n5095);
  and g9121 (n5096, n791, n_4666);
  not g9122 (n_4667, n5096);
  and g9123 (n5097, n795, n_4667);
  not g9124 (n_4668, n5097);
  and g9125 (n5098, n799, n_4668);
  not g9126 (n_4669, n5098);
  and g9127 (n5099, n803, n_4669);
  not g9128 (n_4670, n5099);
  and g9129 (n5100, n807, n_4670);
  not g9130 (n_4671, n5100);
  and g9131 (n5101, n811, n_4671);
  not g9132 (n_4672, n5101);
  and g9133 (n5102, n815, n_4672);
  not g9134 (n_4673, n5102);
  and g9135 (n5103, n819, n_4673);
  not g9136 (n_4674, n5103);
  and g9137 (n5104, n823, n_4674);
  not g9138 (n_4675, n5104);
  and g9139 (n5105, n827, n_4675);
  not g9140 (n_4676, n5105);
  and g9141 (n5106, n831, n_4676);
  not g9142 (n_4677, n5106);
  and g9143 (n5107, n835, n_4677);
  and g9144 (n5108, \req[45] , n_683);
  not g9145 (n_4678, n5107);
  and g9146 (\grant[45] , n_4678, n5108);
  not g9147 (n_4679, n1179);
  and g9148 (n5110, n846, n_4679);
  not g9149 (n_4680, n5110);
  and g9150 (n5111, n851, n_4680);
  not g9151 (n_4681, n5111);
  and g9152 (n5112, n855, n_4681);
  not g9153 (n_4682, n5112);
  and g9154 (n5113, n859, n_4682);
  not g9155 (n_4683, n5113);
  and g9156 (n5114, n863, n_4683);
  not g9157 (n_4684, n5114);
  and g9158 (n5115, n867, n_4684);
  not g9159 (n_4685, n5115);
  and g9160 (n5116, n871, n_4685);
  not g9161 (n_4686, n5116);
  and g9162 (n5117, n875, n_4686);
  not g9163 (n_4687, n5117);
  and g9164 (n5118, n879, n_4687);
  not g9165 (n_4688, n5118);
  and g9166 (n5119, n883, n_4688);
  not g9167 (n_4689, n5119);
  and g9168 (n5120, n887, n_4689);
  not g9169 (n_4690, n5120);
  and g9170 (n5121, n891, n_4690);
  not g9171 (n_4691, n5121);
  and g9172 (n5122, n895, n_4691);
  not g9173 (n_4692, n5122);
  and g9174 (n5123, n899, n_4692);
  not g9175 (n_4693, n5123);
  and g9176 (n5124, n903, n_4693);
  not g9177 (n_4694, n5124);
  and g9178 (n5125, n907, n_4694);
  not g9179 (n_4695, n5125);
  and g9180 (n5126, n911, n_4695);
  not g9181 (n_4696, n5126);
  and g9182 (n5127, n915, n_4696);
  not g9183 (n_4697, n5127);
  and g9184 (n5128, n919, n_4697);
  not g9185 (n_4698, n5128);
  and g9186 (n5129, n923, n_4698);
  not g9187 (n_4699, n5129);
  and g9188 (n5130, n927, n_4699);
  not g9189 (n_4700, n5130);
  and g9190 (n5131, n931, n_4700);
  not g9191 (n_4701, n5131);
  and g9192 (n5132, n935, n_4701);
  not g9193 (n_4702, n5132);
  and g9194 (n5133, n939, n_4702);
  not g9195 (n_4703, n5133);
  and g9196 (n5134, n943, n_4703);
  not g9197 (n_4704, n5134);
  and g9198 (n5135, n947, n_4704);
  not g9199 (n_4705, n5135);
  and g9200 (n5136, n951, n_4705);
  not g9201 (n_4706, n5136);
  and g9202 (n5137, n955, n_4706);
  not g9203 (n_4707, n5137);
  and g9204 (n5138, n959, n_4707);
  not g9205 (n_4708, n5138);
  and g9206 (n5139, n963, n_4708);
  not g9207 (n_4709, n5139);
  and g9208 (n5140, n967, n_4709);
  not g9209 (n_4710, n5140);
  and g9210 (n5141, n971, n_4710);
  not g9211 (n_4711, n5141);
  and g9212 (n5142, n975, n_4711);
  not g9213 (n_4712, n5142);
  and g9214 (n5143, n979, n_4712);
  not g9215 (n_4713, n5143);
  and g9216 (n5144, n983, n_4713);
  not g9217 (n_4714, n5144);
  and g9218 (n5145, n987, n_4714);
  not g9219 (n_4715, n5145);
  and g9220 (n5146, n991, n_4715);
  not g9221 (n_4716, n5146);
  and g9222 (n5147, n995, n_4716);
  not g9223 (n_4717, n5147);
  and g9224 (n5148, n999, n_4717);
  not g9225 (n_4718, n5148);
  and g9226 (n5149, n1003, n_4718);
  not g9227 (n_4719, n5149);
  and g9228 (n5150, n1007, n_4719);
  not g9229 (n_4720, n5150);
  and g9230 (n5151, n1011, n_4720);
  not g9231 (n_4721, n5151);
  and g9232 (n5152, n1015, n_4721);
  not g9233 (n_4722, n5152);
  and g9234 (n5153, n1019, n_4722);
  not g9235 (n_4723, n5153);
  and g9236 (n5154, n1023, n_4723);
  not g9237 (n_4724, n5154);
  and g9238 (n5155, n1027, n_4724);
  not g9239 (n_4725, n5155);
  and g9240 (n5156, n1031, n_4725);
  not g9241 (n_4726, n5156);
  and g9242 (n5157, n1035, n_4726);
  not g9243 (n_4727, n5157);
  and g9244 (n5158, n1039, n_4727);
  not g9245 (n_4728, n5158);
  and g9246 (n5159, n1043, n_4728);
  not g9247 (n_4729, n5159);
  and g9248 (n5160, n1047, n_4729);
  not g9249 (n_4730, n5160);
  and g9250 (n5161, n1051, n_4730);
  not g9251 (n_4731, n5161);
  and g9252 (n5162, n1055, n_4731);
  not g9253 (n_4732, n5162);
  and g9254 (n5163, n1059, n_4732);
  not g9255 (n_4733, n5163);
  and g9256 (n5164, n1574, n_4733);
  not g9257 (n_4734, n5164);
  and g9258 (n5165, n1576, n_4734);
  not g9259 (n_4735, n5165);
  and g9260 (n5166, n1837, n_4735);
  not g9261 (n_4736, n5166);
  and g9262 (n5167, n1068, n_4736);
  not g9263 (n_4737, n5167);
  and g9264 (n5168, n1072, n_4737);
  not g9265 (n_4738, n5168);
  and g9266 (n5169, n1076, n_4738);
  not g9267 (n_4739, n5169);
  and g9268 (n5170, n1080, n_4739);
  not g9269 (n_4740, n5170);
  and g9270 (n5171, n1084, n_4740);
  not g9271 (n_4741, n5171);
  and g9272 (n5172, n1088, n_4741);
  not g9273 (n_4742, n5172);
  and g9274 (n5173, n1092, n_4742);
  not g9275 (n_4743, n5173);
  and g9276 (n5174, n1096, n_4743);
  not g9277 (n_4744, n5174);
  and g9278 (n5175, n1100, n_4744);
  not g9279 (n_4745, n5175);
  and g9280 (n5176, n1104, n_4745);
  not g9281 (n_4746, n5176);
  and g9282 (n5177, n1108, n_4746);
  not g9283 (n_4747, n5177);
  and g9284 (n5178, n1112, n_4747);
  not g9285 (n_4748, n5178);
  and g9286 (n5179, n1116, n_4748);
  not g9287 (n_4749, n5179);
  and g9288 (n5180, n1120, n_4749);
  not g9289 (n_4750, n5180);
  and g9290 (n5181, n1124, n_4750);
  not g9291 (n_4751, n5181);
  and g9292 (n5182, n1128, n_4751);
  not g9293 (n_4752, n5182);
  and g9294 (n5183, n1132, n_4752);
  not g9295 (n_4753, n5183);
  and g9296 (n5184, n1136, n_4753);
  not g9297 (n_4754, n5184);
  and g9298 (n5185, n1140, n_4754);
  not g9299 (n_4755, n5185);
  and g9300 (n5186, n1144, n_4755);
  not g9301 (n_4756, n5186);
  and g9302 (n5187, n1148, n_4756);
  not g9303 (n_4757, n5187);
  and g9304 (n5188, n1152, n_4757);
  not g9305 (n_4758, n5188);
  and g9306 (n5189, n1156, n_4758);
  not g9307 (n_4759, n5189);
  and g9308 (n5190, n1160, n_4759);
  not g9309 (n_4760, n5190);
  and g9310 (n5191, n1164, n_4760);
  not g9311 (n_4761, n5191);
  and g9312 (n5192, n1168, n_4761);
  not g9313 (n_4762, n5192);
  and g9314 (n5193, n1172, n_4762);
  and g9315 (n5194, \req[46] , n_907);
  not g9316 (n_4763, n5193);
  and g9317 (\grant[46] , n_4763, n5194);
  not g9318 (n_4764, n511);
  and g9319 (n5196, n_4764, n1183);
  not g9320 (n_4765, n5196);
  and g9321 (n5197, n1188, n_4765);
  not g9322 (n_4766, n5197);
  and g9323 (n5198, n1192, n_4766);
  not g9324 (n_4767, n5198);
  and g9325 (n5199, n1196, n_4767);
  not g9326 (n_4768, n5199);
  and g9327 (n5200, n1200, n_4768);
  not g9328 (n_4769, n5200);
  and g9329 (n5201, n1204, n_4769);
  not g9330 (n_4770, n5201);
  and g9331 (n5202, n1208, n_4770);
  not g9332 (n_4771, n5202);
  and g9333 (n5203, n1212, n_4771);
  not g9334 (n_4772, n5203);
  and g9335 (n5204, n1216, n_4772);
  not g9336 (n_4773, n5204);
  and g9337 (n5205, n1220, n_4773);
  not g9338 (n_4774, n5205);
  and g9339 (n5206, n1224, n_4774);
  not g9340 (n_4775, n5206);
  and g9341 (n5207, n1228, n_4775);
  not g9342 (n_4776, n5207);
  and g9343 (n5208, n1232, n_4776);
  not g9344 (n_4777, n5208);
  and g9345 (n5209, n1236, n_4777);
  not g9346 (n_4778, n5209);
  and g9347 (n5210, n1240, n_4778);
  not g9348 (n_4779, n5210);
  and g9349 (n5211, n1244, n_4779);
  not g9350 (n_4780, n5211);
  and g9351 (n5212, n1248, n_4780);
  not g9352 (n_4781, n5212);
  and g9353 (n5213, n1252, n_4781);
  not g9354 (n_4782, n5213);
  and g9355 (n5214, n1256, n_4782);
  not g9356 (n_4783, n5214);
  and g9357 (n5215, n1260, n_4783);
  not g9358 (n_4784, n5215);
  and g9359 (n5216, n1264, n_4784);
  not g9360 (n_4785, n5216);
  and g9361 (n5217, n1268, n_4785);
  not g9362 (n_4786, n5217);
  and g9363 (n5218, n1272, n_4786);
  not g9364 (n_4787, n5218);
  and g9365 (n5219, n1276, n_4787);
  not g9366 (n_4788, n5219);
  and g9367 (n5220, n1280, n_4788);
  not g9368 (n_4789, n5220);
  and g9369 (n5221, n1284, n_4789);
  not g9370 (n_4790, n5221);
  and g9371 (n5222, n1288, n_4790);
  not g9372 (n_4791, n5222);
  and g9373 (n5223, n1292, n_4791);
  not g9374 (n_4792, n5223);
  and g9375 (n5224, n1296, n_4792);
  not g9376 (n_4793, n5224);
  and g9377 (n5225, n1300, n_4793);
  not g9378 (n_4794, n5225);
  and g9379 (n5226, n1304, n_4794);
  not g9380 (n_4795, n5226);
  and g9381 (n5227, n1308, n_4795);
  not g9382 (n_4796, n5227);
  and g9383 (n5228, n1312, n_4796);
  not g9384 (n_4797, n5228);
  and g9385 (n5229, n1316, n_4797);
  not g9386 (n_4798, n5229);
  and g9387 (n5230, n1320, n_4798);
  not g9388 (n_4799, n5230);
  and g9389 (n5231, n1324, n_4799);
  not g9390 (n_4800, n5231);
  and g9391 (n5232, n1328, n_4800);
  not g9392 (n_4801, n5232);
  and g9393 (n5233, n1332, n_4801);
  not g9394 (n_4802, n5233);
  and g9395 (n5234, n1336, n_4802);
  not g9396 (n_4803, n5234);
  and g9397 (n5235, n1340, n_4803);
  not g9398 (n_4804, n5235);
  and g9399 (n5236, n1344, n_4804);
  not g9400 (n_4805, n5236);
  and g9401 (n5237, n1348, n_4805);
  not g9402 (n_4806, n5237);
  and g9403 (n5238, n1352, n_4806);
  not g9404 (n_4807, n5238);
  and g9405 (n5239, n1356, n_4807);
  not g9406 (n_4808, n5239);
  and g9407 (n5240, n1360, n_4808);
  not g9408 (n_4809, n5240);
  and g9409 (n5241, n1364, n_4809);
  not g9410 (n_4810, n5241);
  and g9411 (n5242, n1368, n_4810);
  not g9412 (n_4811, n5242);
  and g9413 (n5243, n1372, n_4811);
  not g9414 (n_4812, n5243);
  and g9415 (n5244, n1376, n_4812);
  not g9416 (n_4813, n5244);
  and g9417 (n5245, n1380, n_4813);
  not g9418 (n_4814, n5245);
  and g9419 (n5246, n1384, n_4814);
  not g9420 (n_4815, n5246);
  and g9421 (n5247, n1388, n_4815);
  not g9422 (n_4816, n5247);
  and g9423 (n5248, n1392, n_4816);
  not g9424 (n_4817, n5248);
  and g9425 (n5249, n1396, n_4817);
  not g9426 (n_4818, n5249);
  and g9427 (n5250, n1663, n_4818);
  not g9428 (n_4819, n5250);
  and g9429 (n5251, n392, n_4819);
  not g9430 (n_4820, n5251);
  and g9431 (n5252, n396, n_4820);
  not g9432 (n_4821, n5252);
  and g9433 (n5253, n400, n_4821);
  not g9434 (n_4822, n5253);
  and g9435 (n5254, n404, n_4822);
  not g9436 (n_4823, n5254);
  and g9437 (n5255, n408, n_4823);
  not g9438 (n_4824, n5255);
  and g9439 (n5256, n412, n_4824);
  not g9440 (n_4825, n5256);
  and g9441 (n5257, n416, n_4825);
  not g9442 (n_4826, n5257);
  and g9443 (n5258, n420, n_4826);
  not g9444 (n_4827, n5258);
  and g9445 (n5259, n424, n_4827);
  not g9446 (n_4828, n5259);
  and g9447 (n5260, n428, n_4828);
  not g9448 (n_4829, n5260);
  and g9449 (n5261, n432, n_4829);
  not g9450 (n_4830, n5261);
  and g9451 (n5262, n436, n_4830);
  not g9452 (n_4831, n5262);
  and g9453 (n5263, n440, n_4831);
  not g9454 (n_4832, n5263);
  and g9455 (n5264, n444, n_4832);
  not g9456 (n_4833, n5264);
  and g9457 (n5265, n448, n_4833);
  not g9458 (n_4834, n5265);
  and g9459 (n5266, n452, n_4834);
  not g9460 (n_4835, n5266);
  and g9461 (n5267, n456, n_4835);
  not g9462 (n_4836, n5267);
  and g9463 (n5268, n460, n_4836);
  not g9464 (n_4837, n5268);
  and g9465 (n5269, n464, n_4837);
  not g9466 (n_4838, n5269);
  and g9467 (n5270, n468, n_4838);
  not g9468 (n_4839, n5270);
  and g9469 (n5271, n472, n_4839);
  not g9470 (n_4840, n5271);
  and g9471 (n5272, n476, n_4840);
  not g9472 (n_4841, n5272);
  and g9473 (n5273, n480, n_4841);
  not g9474 (n_4842, n5273);
  and g9475 (n5274, n484, n_4842);
  not g9476 (n_4843, n5274);
  and g9477 (n5275, n488, n_4843);
  not g9478 (n_4844, n5275);
  and g9479 (n5276, n492, n_4844);
  not g9480 (n_4845, n5276);
  and g9481 (n5277, n496, n_4845);
  not g9482 (n_4846, n5277);
  and g9483 (n5278, n500, n_4846);
  not g9484 (n_4847, n5278);
  and g9485 (n5279, n504, n_4847);
  and g9486 (n5280, \req[47] , n_220);
  not g9487 (n_4848, n5279);
  and g9488 (\grant[47] , n_4848, n5280);
  not g9489 (n_4849, n850);
  and g9490 (n5282, n515, n_4849);
  not g9491 (n_4850, n5282);
  and g9492 (n5283, n520, n_4850);
  not g9493 (n_4851, n5283);
  and g9494 (n5284, n524, n_4851);
  not g9495 (n_4852, n5284);
  and g9496 (n5285, n528, n_4852);
  not g9497 (n_4853, n5285);
  and g9498 (n5286, n532, n_4853);
  not g9499 (n_4854, n5286);
  and g9500 (n5287, n536, n_4854);
  not g9501 (n_4855, n5287);
  and g9502 (n5288, n540, n_4855);
  not g9503 (n_4856, n5288);
  and g9504 (n5289, n544, n_4856);
  not g9505 (n_4857, n5289);
  and g9506 (n5290, n548, n_4857);
  not g9507 (n_4858, n5290);
  and g9508 (n5291, n552, n_4858);
  not g9509 (n_4859, n5291);
  and g9510 (n5292, n556, n_4859);
  not g9511 (n_4860, n5292);
  and g9512 (n5293, n560, n_4860);
  not g9513 (n_4861, n5293);
  and g9514 (n5294, n564, n_4861);
  not g9515 (n_4862, n5294);
  and g9516 (n5295, n568, n_4862);
  not g9517 (n_4863, n5295);
  and g9518 (n5296, n572, n_4863);
  not g9519 (n_4864, n5296);
  and g9520 (n5297, n576, n_4864);
  not g9521 (n_4865, n5297);
  and g9522 (n5298, n580, n_4865);
  not g9523 (n_4866, n5298);
  and g9524 (n5299, n584, n_4866);
  not g9525 (n_4867, n5299);
  and g9526 (n5300, n588, n_4867);
  not g9527 (n_4868, n5300);
  and g9528 (n5301, n592, n_4868);
  not g9529 (n_4869, n5301);
  and g9530 (n5302, n596, n_4869);
  not g9531 (n_4870, n5302);
  and g9532 (n5303, n600, n_4870);
  not g9533 (n_4871, n5303);
  and g9534 (n5304, n604, n_4871);
  not g9535 (n_4872, n5304);
  and g9536 (n5305, n608, n_4872);
  not g9537 (n_4873, n5305);
  and g9538 (n5306, n612, n_4873);
  not g9539 (n_4874, n5306);
  and g9540 (n5307, n616, n_4874);
  not g9541 (n_4875, n5307);
  and g9542 (n5308, n620, n_4875);
  not g9543 (n_4876, n5308);
  and g9544 (n5309, n624, n_4876);
  not g9545 (n_4877, n5309);
  and g9546 (n5310, n628, n_4877);
  not g9547 (n_4878, n5310);
  and g9548 (n5311, n632, n_4878);
  not g9549 (n_4879, n5311);
  and g9550 (n5312, n636, n_4879);
  not g9551 (n_4880, n5312);
  and g9552 (n5313, n640, n_4880);
  not g9553 (n_4881, n5313);
  and g9554 (n5314, n644, n_4881);
  not g9555 (n_4882, n5314);
  and g9556 (n5315, n648, n_4882);
  not g9557 (n_4883, n5315);
  and g9558 (n5316, n652, n_4883);
  not g9559 (n_4884, n5316);
  and g9560 (n5317, n656, n_4884);
  not g9561 (n_4885, n5317);
  and g9562 (n5318, n660, n_4885);
  not g9563 (n_4886, n5318);
  and g9564 (n5319, n664, n_4886);
  not g9565 (n_4887, n5319);
  and g9566 (n5320, n668, n_4887);
  not g9567 (n_4888, n5320);
  and g9568 (n5321, n672, n_4888);
  not g9569 (n_4889, n5321);
  and g9570 (n5322, n676, n_4889);
  not g9571 (n_4890, n5322);
  and g9572 (n5323, n680, n_4890);
  not g9573 (n_4891, n5323);
  and g9574 (n5324, n684, n_4891);
  not g9575 (n_4892, n5324);
  and g9576 (n5325, n688, n_4892);
  not g9577 (n_4893, n5325);
  and g9578 (n5326, n692, n_4893);
  not g9579 (n_4894, n5326);
  and g9580 (n5327, n696, n_4894);
  not g9581 (n_4895, n5327);
  and g9582 (n5328, n700, n_4895);
  not g9583 (n_4896, n5328);
  and g9584 (n5329, n704, n_4896);
  not g9585 (n_4897, n5329);
  and g9586 (n5330, n708, n_4897);
  not g9587 (n_4898, n5330);
  and g9588 (n5331, n712, n_4898);
  not g9589 (n_4899, n5331);
  and g9590 (n5332, n716, n_4899);
  not g9591 (n_4900, n5332);
  and g9592 (n5333, n720, n_4900);
  not g9593 (n_4901, n5333);
  and g9594 (n5334, n1484, n_4901);
  not g9595 (n_4902, n5334);
  and g9596 (n5335, n1486, n_4902);
  not g9597 (n_4903, n5335);
  and g9598 (n5336, n1750, n_4903);
  not g9599 (n_4904, n5336);
  and g9600 (n5337, n731, n_4904);
  not g9601 (n_4905, n5337);
  and g9602 (n5338, n735, n_4905);
  not g9603 (n_4906, n5338);
  and g9604 (n5339, n739, n_4906);
  not g9605 (n_4907, n5339);
  and g9606 (n5340, n743, n_4907);
  not g9607 (n_4908, n5340);
  and g9608 (n5341, n747, n_4908);
  not g9609 (n_4909, n5341);
  and g9610 (n5342, n751, n_4909);
  not g9611 (n_4910, n5342);
  and g9612 (n5343, n755, n_4910);
  not g9613 (n_4911, n5343);
  and g9614 (n5344, n759, n_4911);
  not g9615 (n_4912, n5344);
  and g9616 (n5345, n763, n_4912);
  not g9617 (n_4913, n5345);
  and g9618 (n5346, n767, n_4913);
  not g9619 (n_4914, n5346);
  and g9620 (n5347, n771, n_4914);
  not g9621 (n_4915, n5347);
  and g9622 (n5348, n775, n_4915);
  not g9623 (n_4916, n5348);
  and g9624 (n5349, n779, n_4916);
  not g9625 (n_4917, n5349);
  and g9626 (n5350, n783, n_4917);
  not g9627 (n_4918, n5350);
  and g9628 (n5351, n787, n_4918);
  not g9629 (n_4919, n5351);
  and g9630 (n5352, n791, n_4919);
  not g9631 (n_4920, n5352);
  and g9632 (n5353, n795, n_4920);
  not g9633 (n_4921, n5353);
  and g9634 (n5354, n799, n_4921);
  not g9635 (n_4922, n5354);
  and g9636 (n5355, n803, n_4922);
  not g9637 (n_4923, n5355);
  and g9638 (n5356, n807, n_4923);
  not g9639 (n_4924, n5356);
  and g9640 (n5357, n811, n_4924);
  not g9641 (n_4925, n5357);
  and g9642 (n5358, n815, n_4925);
  not g9643 (n_4926, n5358);
  and g9644 (n5359, n819, n_4926);
  not g9645 (n_4927, n5359);
  and g9646 (n5360, n823, n_4927);
  not g9647 (n_4928, n5360);
  and g9648 (n5361, n827, n_4928);
  not g9649 (n_4929, n5361);
  and g9650 (n5362, n831, n_4929);
  not g9651 (n_4930, n5362);
  and g9652 (n5363, n835, n_4930);
  not g9653 (n_4931, n5363);
  and g9654 (n5364, n839, n_4931);
  not g9655 (n_4932, n5364);
  and g9656 (n5365, n843, n_4932);
  and g9657 (n5366, \req[48] , n_689);
  not g9658 (n_4933, n5365);
  and g9659 (\grant[48] , n_4933, n5366);
  not g9660 (n_4934, n1187);
  and g9661 (n5368, n854, n_4934);
  not g9662 (n_4935, n5368);
  and g9663 (n5369, n859, n_4935);
  not g9664 (n_4936, n5369);
  and g9665 (n5370, n863, n_4936);
  not g9666 (n_4937, n5370);
  and g9667 (n5371, n867, n_4937);
  not g9668 (n_4938, n5371);
  and g9669 (n5372, n871, n_4938);
  not g9670 (n_4939, n5372);
  and g9671 (n5373, n875, n_4939);
  not g9672 (n_4940, n5373);
  and g9673 (n5374, n879, n_4940);
  not g9674 (n_4941, n5374);
  and g9675 (n5375, n883, n_4941);
  not g9676 (n_4942, n5375);
  and g9677 (n5376, n887, n_4942);
  not g9678 (n_4943, n5376);
  and g9679 (n5377, n891, n_4943);
  not g9680 (n_4944, n5377);
  and g9681 (n5378, n895, n_4944);
  not g9682 (n_4945, n5378);
  and g9683 (n5379, n899, n_4945);
  not g9684 (n_4946, n5379);
  and g9685 (n5380, n903, n_4946);
  not g9686 (n_4947, n5380);
  and g9687 (n5381, n907, n_4947);
  not g9688 (n_4948, n5381);
  and g9689 (n5382, n911, n_4948);
  not g9690 (n_4949, n5382);
  and g9691 (n5383, n915, n_4949);
  not g9692 (n_4950, n5383);
  and g9693 (n5384, n919, n_4950);
  not g9694 (n_4951, n5384);
  and g9695 (n5385, n923, n_4951);
  not g9696 (n_4952, n5385);
  and g9697 (n5386, n927, n_4952);
  not g9698 (n_4953, n5386);
  and g9699 (n5387, n931, n_4953);
  not g9700 (n_4954, n5387);
  and g9701 (n5388, n935, n_4954);
  not g9702 (n_4955, n5388);
  and g9703 (n5389, n939, n_4955);
  not g9704 (n_4956, n5389);
  and g9705 (n5390, n943, n_4956);
  not g9706 (n_4957, n5390);
  and g9707 (n5391, n947, n_4957);
  not g9708 (n_4958, n5391);
  and g9709 (n5392, n951, n_4958);
  not g9710 (n_4959, n5392);
  and g9711 (n5393, n955, n_4959);
  not g9712 (n_4960, n5393);
  and g9713 (n5394, n959, n_4960);
  not g9714 (n_4961, n5394);
  and g9715 (n5395, n963, n_4961);
  not g9716 (n_4962, n5395);
  and g9717 (n5396, n967, n_4962);
  not g9718 (n_4963, n5396);
  and g9719 (n5397, n971, n_4963);
  not g9720 (n_4964, n5397);
  and g9721 (n5398, n975, n_4964);
  not g9722 (n_4965, n5398);
  and g9723 (n5399, n979, n_4965);
  not g9724 (n_4966, n5399);
  and g9725 (n5400, n983, n_4966);
  not g9726 (n_4967, n5400);
  and g9727 (n5401, n987, n_4967);
  not g9728 (n_4968, n5401);
  and g9729 (n5402, n991, n_4968);
  not g9730 (n_4969, n5402);
  and g9731 (n5403, n995, n_4969);
  not g9732 (n_4970, n5403);
  and g9733 (n5404, n999, n_4970);
  not g9734 (n_4971, n5404);
  and g9735 (n5405, n1003, n_4971);
  not g9736 (n_4972, n5405);
  and g9737 (n5406, n1007, n_4972);
  not g9738 (n_4973, n5406);
  and g9739 (n5407, n1011, n_4973);
  not g9740 (n_4974, n5407);
  and g9741 (n5408, n1015, n_4974);
  not g9742 (n_4975, n5408);
  and g9743 (n5409, n1019, n_4975);
  not g9744 (n_4976, n5409);
  and g9745 (n5410, n1023, n_4976);
  not g9746 (n_4977, n5410);
  and g9747 (n5411, n1027, n_4977);
  not g9748 (n_4978, n5411);
  and g9749 (n5412, n1031, n_4978);
  not g9750 (n_4979, n5412);
  and g9751 (n5413, n1035, n_4979);
  not g9752 (n_4980, n5413);
  and g9753 (n5414, n1039, n_4980);
  not g9754 (n_4981, n5414);
  and g9755 (n5415, n1043, n_4981);
  not g9756 (n_4982, n5415);
  and g9757 (n5416, n1047, n_4982);
  not g9758 (n_4983, n5416);
  and g9759 (n5417, n1051, n_4983);
  not g9760 (n_4984, n5417);
  and g9761 (n5418, n1055, n_4984);
  not g9762 (n_4985, n5418);
  and g9763 (n5419, n1059, n_4985);
  not g9764 (n_4986, n5419);
  and g9765 (n5420, n1574, n_4986);
  not g9766 (n_4987, n5420);
  and g9767 (n5421, n1576, n_4987);
  not g9768 (n_4988, n5421);
  and g9769 (n5422, n1837, n_4988);
  not g9770 (n_4989, n5422);
  and g9771 (n5423, n1068, n_4989);
  not g9772 (n_4990, n5423);
  and g9773 (n5424, n1072, n_4990);
  not g9774 (n_4991, n5424);
  and g9775 (n5425, n1076, n_4991);
  not g9776 (n_4992, n5425);
  and g9777 (n5426, n1080, n_4992);
  not g9778 (n_4993, n5426);
  and g9779 (n5427, n1084, n_4993);
  not g9780 (n_4994, n5427);
  and g9781 (n5428, n1088, n_4994);
  not g9782 (n_4995, n5428);
  and g9783 (n5429, n1092, n_4995);
  not g9784 (n_4996, n5429);
  and g9785 (n5430, n1096, n_4996);
  not g9786 (n_4997, n5430);
  and g9787 (n5431, n1100, n_4997);
  not g9788 (n_4998, n5431);
  and g9789 (n5432, n1104, n_4998);
  not g9790 (n_4999, n5432);
  and g9791 (n5433, n1108, n_4999);
  not g9792 (n_5000, n5433);
  and g9793 (n5434, n1112, n_5000);
  not g9794 (n_5001, n5434);
  and g9795 (n5435, n1116, n_5001);
  not g9796 (n_5002, n5435);
  and g9797 (n5436, n1120, n_5002);
  not g9798 (n_5003, n5436);
  and g9799 (n5437, n1124, n_5003);
  not g9800 (n_5004, n5437);
  and g9801 (n5438, n1128, n_5004);
  not g9802 (n_5005, n5438);
  and g9803 (n5439, n1132, n_5005);
  not g9804 (n_5006, n5439);
  and g9805 (n5440, n1136, n_5006);
  not g9806 (n_5007, n5440);
  and g9807 (n5441, n1140, n_5007);
  not g9808 (n_5008, n5441);
  and g9809 (n5442, n1144, n_5008);
  not g9810 (n_5009, n5442);
  and g9811 (n5443, n1148, n_5009);
  not g9812 (n_5010, n5443);
  and g9813 (n5444, n1152, n_5010);
  not g9814 (n_5011, n5444);
  and g9815 (n5445, n1156, n_5011);
  not g9816 (n_5012, n5445);
  and g9817 (n5446, n1160, n_5012);
  not g9818 (n_5013, n5446);
  and g9819 (n5447, n1164, n_5013);
  not g9820 (n_5014, n5447);
  and g9821 (n5448, n1168, n_5014);
  not g9822 (n_5015, n5448);
  and g9823 (n5449, n1172, n_5015);
  not g9824 (n_5016, n5449);
  and g9825 (n5450, n1176, n_5016);
  not g9826 (n_5017, n5450);
  and g9827 (n5451, n1180, n_5017);
  and g9828 (n5452, \req[49] , n_911);
  not g9829 (n_5018, n5451);
  and g9830 (\grant[49] , n_5018, n5452);
  not g9831 (n_5019, n519);
  and g9832 (n5454, n_5019, n1191);
  not g9833 (n_5020, n5454);
  and g9834 (n5455, n1196, n_5020);
  not g9835 (n_5021, n5455);
  and g9836 (n5456, n1200, n_5021);
  not g9837 (n_5022, n5456);
  and g9838 (n5457, n1204, n_5022);
  not g9839 (n_5023, n5457);
  and g9840 (n5458, n1208, n_5023);
  not g9841 (n_5024, n5458);
  and g9842 (n5459, n1212, n_5024);
  not g9843 (n_5025, n5459);
  and g9844 (n5460, n1216, n_5025);
  not g9845 (n_5026, n5460);
  and g9846 (n5461, n1220, n_5026);
  not g9847 (n_5027, n5461);
  and g9848 (n5462, n1224, n_5027);
  not g9849 (n_5028, n5462);
  and g9850 (n5463, n1228, n_5028);
  not g9851 (n_5029, n5463);
  and g9852 (n5464, n1232, n_5029);
  not g9853 (n_5030, n5464);
  and g9854 (n5465, n1236, n_5030);
  not g9855 (n_5031, n5465);
  and g9856 (n5466, n1240, n_5031);
  not g9857 (n_5032, n5466);
  and g9858 (n5467, n1244, n_5032);
  not g9859 (n_5033, n5467);
  and g9860 (n5468, n1248, n_5033);
  not g9861 (n_5034, n5468);
  and g9862 (n5469, n1252, n_5034);
  not g9863 (n_5035, n5469);
  and g9864 (n5470, n1256, n_5035);
  not g9865 (n_5036, n5470);
  and g9866 (n5471, n1260, n_5036);
  not g9867 (n_5037, n5471);
  and g9868 (n5472, n1264, n_5037);
  not g9869 (n_5038, n5472);
  and g9870 (n5473, n1268, n_5038);
  not g9871 (n_5039, n5473);
  and g9872 (n5474, n1272, n_5039);
  not g9873 (n_5040, n5474);
  and g9874 (n5475, n1276, n_5040);
  not g9875 (n_5041, n5475);
  and g9876 (n5476, n1280, n_5041);
  not g9877 (n_5042, n5476);
  and g9878 (n5477, n1284, n_5042);
  not g9879 (n_5043, n5477);
  and g9880 (n5478, n1288, n_5043);
  not g9881 (n_5044, n5478);
  and g9882 (n5479, n1292, n_5044);
  not g9883 (n_5045, n5479);
  and g9884 (n5480, n1296, n_5045);
  not g9885 (n_5046, n5480);
  and g9886 (n5481, n1300, n_5046);
  not g9887 (n_5047, n5481);
  and g9888 (n5482, n1304, n_5047);
  not g9889 (n_5048, n5482);
  and g9890 (n5483, n1308, n_5048);
  not g9891 (n_5049, n5483);
  and g9892 (n5484, n1312, n_5049);
  not g9893 (n_5050, n5484);
  and g9894 (n5485, n1316, n_5050);
  not g9895 (n_5051, n5485);
  and g9896 (n5486, n1320, n_5051);
  not g9897 (n_5052, n5486);
  and g9898 (n5487, n1324, n_5052);
  not g9899 (n_5053, n5487);
  and g9900 (n5488, n1328, n_5053);
  not g9901 (n_5054, n5488);
  and g9902 (n5489, n1332, n_5054);
  not g9903 (n_5055, n5489);
  and g9904 (n5490, n1336, n_5055);
  not g9905 (n_5056, n5490);
  and g9906 (n5491, n1340, n_5056);
  not g9907 (n_5057, n5491);
  and g9908 (n5492, n1344, n_5057);
  not g9909 (n_5058, n5492);
  and g9910 (n5493, n1348, n_5058);
  not g9911 (n_5059, n5493);
  and g9912 (n5494, n1352, n_5059);
  not g9913 (n_5060, n5494);
  and g9914 (n5495, n1356, n_5060);
  not g9915 (n_5061, n5495);
  and g9916 (n5496, n1360, n_5061);
  not g9917 (n_5062, n5496);
  and g9918 (n5497, n1364, n_5062);
  not g9919 (n_5063, n5497);
  and g9920 (n5498, n1368, n_5063);
  not g9921 (n_5064, n5498);
  and g9922 (n5499, n1372, n_5064);
  not g9923 (n_5065, n5499);
  and g9924 (n5500, n1376, n_5065);
  not g9925 (n_5066, n5500);
  and g9926 (n5501, n1380, n_5066);
  not g9927 (n_5067, n5501);
  and g9928 (n5502, n1384, n_5067);
  not g9929 (n_5068, n5502);
  and g9930 (n5503, n1388, n_5068);
  not g9931 (n_5069, n5503);
  and g9932 (n5504, n1392, n_5069);
  not g9933 (n_5070, n5504);
  and g9934 (n5505, n1396, n_5070);
  not g9935 (n_5071, n5505);
  and g9936 (n5506, n1663, n_5071);
  not g9937 (n_5072, n5506);
  and g9938 (n5507, n392, n_5072);
  not g9939 (n_5073, n5507);
  and g9940 (n5508, n396, n_5073);
  not g9941 (n_5074, n5508);
  and g9942 (n5509, n400, n_5074);
  not g9943 (n_5075, n5509);
  and g9944 (n5510, n404, n_5075);
  not g9945 (n_5076, n5510);
  and g9946 (n5511, n408, n_5076);
  not g9947 (n_5077, n5511);
  and g9948 (n5512, n412, n_5077);
  not g9949 (n_5078, n5512);
  and g9950 (n5513, n416, n_5078);
  not g9951 (n_5079, n5513);
  and g9952 (n5514, n420, n_5079);
  not g9953 (n_5080, n5514);
  and g9954 (n5515, n424, n_5080);
  not g9955 (n_5081, n5515);
  and g9956 (n5516, n428, n_5081);
  not g9957 (n_5082, n5516);
  and g9958 (n5517, n432, n_5082);
  not g9959 (n_5083, n5517);
  and g9960 (n5518, n436, n_5083);
  not g9961 (n_5084, n5518);
  and g9962 (n5519, n440, n_5084);
  not g9963 (n_5085, n5519);
  and g9964 (n5520, n444, n_5085);
  not g9965 (n_5086, n5520);
  and g9966 (n5521, n448, n_5086);
  not g9967 (n_5087, n5521);
  and g9968 (n5522, n452, n_5087);
  not g9969 (n_5088, n5522);
  and g9970 (n5523, n456, n_5088);
  not g9971 (n_5089, n5523);
  and g9972 (n5524, n460, n_5089);
  not g9973 (n_5090, n5524);
  and g9974 (n5525, n464, n_5090);
  not g9975 (n_5091, n5525);
  and g9976 (n5526, n468, n_5091);
  not g9977 (n_5092, n5526);
  and g9978 (n5527, n472, n_5092);
  not g9979 (n_5093, n5527);
  and g9980 (n5528, n476, n_5093);
  not g9981 (n_5094, n5528);
  and g9982 (n5529, n480, n_5094);
  not g9983 (n_5095, n5529);
  and g9984 (n5530, n484, n_5095);
  not g9985 (n_5096, n5530);
  and g9986 (n5531, n488, n_5096);
  not g9987 (n_5097, n5531);
  and g9988 (n5532, n492, n_5097);
  not g9989 (n_5098, n5532);
  and g9990 (n5533, n496, n_5098);
  not g9991 (n_5099, n5533);
  and g9992 (n5534, n500, n_5099);
  not g9993 (n_5100, n5534);
  and g9994 (n5535, n504, n_5100);
  not g9995 (n_5101, n5535);
  and g9996 (n5536, n508, n_5101);
  not g9997 (n_5102, n5536);
  and g9998 (n5537, n512, n_5102);
  and g9999 (n5538, \req[50] , n_234);
  not g10000 (n_5103, n5537);
  and g10001 (\grant[50] , n_5103, n5538);
  not g10002 (n_5104, n858);
  and g10003 (n5540, n523, n_5104);
  not g10004 (n_5105, n5540);
  and g10005 (n5541, n528, n_5105);
  not g10006 (n_5106, n5541);
  and g10007 (n5542, n532, n_5106);
  not g10008 (n_5107, n5542);
  and g10009 (n5543, n536, n_5107);
  not g10010 (n_5108, n5543);
  and g10011 (n5544, n540, n_5108);
  not g10012 (n_5109, n5544);
  and g10013 (n5545, n544, n_5109);
  not g10014 (n_5110, n5545);
  and g10015 (n5546, n548, n_5110);
  not g10016 (n_5111, n5546);
  and g10017 (n5547, n552, n_5111);
  not g10018 (n_5112, n5547);
  and g10019 (n5548, n556, n_5112);
  not g10020 (n_5113, n5548);
  and g10021 (n5549, n560, n_5113);
  not g10022 (n_5114, n5549);
  and g10023 (n5550, n564, n_5114);
  not g10024 (n_5115, n5550);
  and g10025 (n5551, n568, n_5115);
  not g10026 (n_5116, n5551);
  and g10027 (n5552, n572, n_5116);
  not g10028 (n_5117, n5552);
  and g10029 (n5553, n576, n_5117);
  not g10030 (n_5118, n5553);
  and g10031 (n5554, n580, n_5118);
  not g10032 (n_5119, n5554);
  and g10033 (n5555, n584, n_5119);
  not g10034 (n_5120, n5555);
  and g10035 (n5556, n588, n_5120);
  not g10036 (n_5121, n5556);
  and g10037 (n5557, n592, n_5121);
  not g10038 (n_5122, n5557);
  and g10039 (n5558, n596, n_5122);
  not g10040 (n_5123, n5558);
  and g10041 (n5559, n600, n_5123);
  not g10042 (n_5124, n5559);
  and g10043 (n5560, n604, n_5124);
  not g10044 (n_5125, n5560);
  and g10045 (n5561, n608, n_5125);
  not g10046 (n_5126, n5561);
  and g10047 (n5562, n612, n_5126);
  not g10048 (n_5127, n5562);
  and g10049 (n5563, n616, n_5127);
  not g10050 (n_5128, n5563);
  and g10051 (n5564, n620, n_5128);
  not g10052 (n_5129, n5564);
  and g10053 (n5565, n624, n_5129);
  not g10054 (n_5130, n5565);
  and g10055 (n5566, n628, n_5130);
  not g10056 (n_5131, n5566);
  and g10057 (n5567, n632, n_5131);
  not g10058 (n_5132, n5567);
  and g10059 (n5568, n636, n_5132);
  not g10060 (n_5133, n5568);
  and g10061 (n5569, n640, n_5133);
  not g10062 (n_5134, n5569);
  and g10063 (n5570, n644, n_5134);
  not g10064 (n_5135, n5570);
  and g10065 (n5571, n648, n_5135);
  not g10066 (n_5136, n5571);
  and g10067 (n5572, n652, n_5136);
  not g10068 (n_5137, n5572);
  and g10069 (n5573, n656, n_5137);
  not g10070 (n_5138, n5573);
  and g10071 (n5574, n660, n_5138);
  not g10072 (n_5139, n5574);
  and g10073 (n5575, n664, n_5139);
  not g10074 (n_5140, n5575);
  and g10075 (n5576, n668, n_5140);
  not g10076 (n_5141, n5576);
  and g10077 (n5577, n672, n_5141);
  not g10078 (n_5142, n5577);
  and g10079 (n5578, n676, n_5142);
  not g10080 (n_5143, n5578);
  and g10081 (n5579, n680, n_5143);
  not g10082 (n_5144, n5579);
  and g10083 (n5580, n684, n_5144);
  not g10084 (n_5145, n5580);
  and g10085 (n5581, n688, n_5145);
  not g10086 (n_5146, n5581);
  and g10087 (n5582, n692, n_5146);
  not g10088 (n_5147, n5582);
  and g10089 (n5583, n696, n_5147);
  not g10090 (n_5148, n5583);
  and g10091 (n5584, n700, n_5148);
  not g10092 (n_5149, n5584);
  and g10093 (n5585, n704, n_5149);
  not g10094 (n_5150, n5585);
  and g10095 (n5586, n708, n_5150);
  not g10096 (n_5151, n5586);
  and g10097 (n5587, n712, n_5151);
  not g10098 (n_5152, n5587);
  and g10099 (n5588, n716, n_5152);
  not g10100 (n_5153, n5588);
  and g10101 (n5589, n720, n_5153);
  not g10102 (n_5154, n5589);
  and g10103 (n5590, n1484, n_5154);
  not g10104 (n_5155, n5590);
  and g10105 (n5591, n1486, n_5155);
  not g10106 (n_5156, n5591);
  and g10107 (n5592, n1750, n_5156);
  not g10108 (n_5157, n5592);
  and g10109 (n5593, n731, n_5157);
  not g10110 (n_5158, n5593);
  and g10111 (n5594, n735, n_5158);
  not g10112 (n_5159, n5594);
  and g10113 (n5595, n739, n_5159);
  not g10114 (n_5160, n5595);
  and g10115 (n5596, n743, n_5160);
  not g10116 (n_5161, n5596);
  and g10117 (n5597, n747, n_5161);
  not g10118 (n_5162, n5597);
  and g10119 (n5598, n751, n_5162);
  not g10120 (n_5163, n5598);
  and g10121 (n5599, n755, n_5163);
  not g10122 (n_5164, n5599);
  and g10123 (n5600, n759, n_5164);
  not g10124 (n_5165, n5600);
  and g10125 (n5601, n763, n_5165);
  not g10126 (n_5166, n5601);
  and g10127 (n5602, n767, n_5166);
  not g10128 (n_5167, n5602);
  and g10129 (n5603, n771, n_5167);
  not g10130 (n_5168, n5603);
  and g10131 (n5604, n775, n_5168);
  not g10132 (n_5169, n5604);
  and g10133 (n5605, n779, n_5169);
  not g10134 (n_5170, n5605);
  and g10135 (n5606, n783, n_5170);
  not g10136 (n_5171, n5606);
  and g10137 (n5607, n787, n_5171);
  not g10138 (n_5172, n5607);
  and g10139 (n5608, n791, n_5172);
  not g10140 (n_5173, n5608);
  and g10141 (n5609, n795, n_5173);
  not g10142 (n_5174, n5609);
  and g10143 (n5610, n799, n_5174);
  not g10144 (n_5175, n5610);
  and g10145 (n5611, n803, n_5175);
  not g10146 (n_5176, n5611);
  and g10147 (n5612, n807, n_5176);
  not g10148 (n_5177, n5612);
  and g10149 (n5613, n811, n_5177);
  not g10150 (n_5178, n5613);
  and g10151 (n5614, n815, n_5178);
  not g10152 (n_5179, n5614);
  and g10153 (n5615, n819, n_5179);
  not g10154 (n_5180, n5615);
  and g10155 (n5616, n823, n_5180);
  not g10156 (n_5181, n5616);
  and g10157 (n5617, n827, n_5181);
  not g10158 (n_5182, n5617);
  and g10159 (n5618, n831, n_5182);
  not g10160 (n_5183, n5618);
  and g10161 (n5619, n835, n_5183);
  not g10162 (n_5184, n5619);
  and g10163 (n5620, n839, n_5184);
  not g10164 (n_5185, n5620);
  and g10165 (n5621, n843, n_5185);
  not g10166 (n_5186, n5621);
  and g10167 (n5622, n847, n_5186);
  not g10168 (n_5187, n5622);
  and g10169 (n5623, n851, n_5187);
  and g10170 (n5624, \req[51] , n_695);
  not g10171 (n_5188, n5623);
  and g10172 (\grant[51] , n_5188, n5624);
  not g10173 (n_5189, n1195);
  and g10174 (n5626, n862, n_5189);
  not g10175 (n_5190, n5626);
  and g10176 (n5627, n867, n_5190);
  not g10177 (n_5191, n5627);
  and g10178 (n5628, n871, n_5191);
  not g10179 (n_5192, n5628);
  and g10180 (n5629, n875, n_5192);
  not g10181 (n_5193, n5629);
  and g10182 (n5630, n879, n_5193);
  not g10183 (n_5194, n5630);
  and g10184 (n5631, n883, n_5194);
  not g10185 (n_5195, n5631);
  and g10186 (n5632, n887, n_5195);
  not g10187 (n_5196, n5632);
  and g10188 (n5633, n891, n_5196);
  not g10189 (n_5197, n5633);
  and g10190 (n5634, n895, n_5197);
  not g10191 (n_5198, n5634);
  and g10192 (n5635, n899, n_5198);
  not g10193 (n_5199, n5635);
  and g10194 (n5636, n903, n_5199);
  not g10195 (n_5200, n5636);
  and g10196 (n5637, n907, n_5200);
  not g10197 (n_5201, n5637);
  and g10198 (n5638, n911, n_5201);
  not g10199 (n_5202, n5638);
  and g10200 (n5639, n915, n_5202);
  not g10201 (n_5203, n5639);
  and g10202 (n5640, n919, n_5203);
  not g10203 (n_5204, n5640);
  and g10204 (n5641, n923, n_5204);
  not g10205 (n_5205, n5641);
  and g10206 (n5642, n927, n_5205);
  not g10207 (n_5206, n5642);
  and g10208 (n5643, n931, n_5206);
  not g10209 (n_5207, n5643);
  and g10210 (n5644, n935, n_5207);
  not g10211 (n_5208, n5644);
  and g10212 (n5645, n939, n_5208);
  not g10213 (n_5209, n5645);
  and g10214 (n5646, n943, n_5209);
  not g10215 (n_5210, n5646);
  and g10216 (n5647, n947, n_5210);
  not g10217 (n_5211, n5647);
  and g10218 (n5648, n951, n_5211);
  not g10219 (n_5212, n5648);
  and g10220 (n5649, n955, n_5212);
  not g10221 (n_5213, n5649);
  and g10222 (n5650, n959, n_5213);
  not g10223 (n_5214, n5650);
  and g10224 (n5651, n963, n_5214);
  not g10225 (n_5215, n5651);
  and g10226 (n5652, n967, n_5215);
  not g10227 (n_5216, n5652);
  and g10228 (n5653, n971, n_5216);
  not g10229 (n_5217, n5653);
  and g10230 (n5654, n975, n_5217);
  not g10231 (n_5218, n5654);
  and g10232 (n5655, n979, n_5218);
  not g10233 (n_5219, n5655);
  and g10234 (n5656, n983, n_5219);
  not g10235 (n_5220, n5656);
  and g10236 (n5657, n987, n_5220);
  not g10237 (n_5221, n5657);
  and g10238 (n5658, n991, n_5221);
  not g10239 (n_5222, n5658);
  and g10240 (n5659, n995, n_5222);
  not g10241 (n_5223, n5659);
  and g10242 (n5660, n999, n_5223);
  not g10243 (n_5224, n5660);
  and g10244 (n5661, n1003, n_5224);
  not g10245 (n_5225, n5661);
  and g10246 (n5662, n1007, n_5225);
  not g10247 (n_5226, n5662);
  and g10248 (n5663, n1011, n_5226);
  not g10249 (n_5227, n5663);
  and g10250 (n5664, n1015, n_5227);
  not g10251 (n_5228, n5664);
  and g10252 (n5665, n1019, n_5228);
  not g10253 (n_5229, n5665);
  and g10254 (n5666, n1023, n_5229);
  not g10255 (n_5230, n5666);
  and g10256 (n5667, n1027, n_5230);
  not g10257 (n_5231, n5667);
  and g10258 (n5668, n1031, n_5231);
  not g10259 (n_5232, n5668);
  and g10260 (n5669, n1035, n_5232);
  not g10261 (n_5233, n5669);
  and g10262 (n5670, n1039, n_5233);
  not g10263 (n_5234, n5670);
  and g10264 (n5671, n1043, n_5234);
  not g10265 (n_5235, n5671);
  and g10266 (n5672, n1047, n_5235);
  not g10267 (n_5236, n5672);
  and g10268 (n5673, n1051, n_5236);
  not g10269 (n_5237, n5673);
  and g10270 (n5674, n1055, n_5237);
  not g10271 (n_5238, n5674);
  and g10272 (n5675, n1059, n_5238);
  not g10273 (n_5239, n5675);
  and g10274 (n5676, n1574, n_5239);
  not g10275 (n_5240, n5676);
  and g10276 (n5677, n1576, n_5240);
  not g10277 (n_5241, n5677);
  and g10278 (n5678, n1837, n_5241);
  not g10279 (n_5242, n5678);
  and g10280 (n5679, n1068, n_5242);
  not g10281 (n_5243, n5679);
  and g10282 (n5680, n1072, n_5243);
  not g10283 (n_5244, n5680);
  and g10284 (n5681, n1076, n_5244);
  not g10285 (n_5245, n5681);
  and g10286 (n5682, n1080, n_5245);
  not g10287 (n_5246, n5682);
  and g10288 (n5683, n1084, n_5246);
  not g10289 (n_5247, n5683);
  and g10290 (n5684, n1088, n_5247);
  not g10291 (n_5248, n5684);
  and g10292 (n5685, n1092, n_5248);
  not g10293 (n_5249, n5685);
  and g10294 (n5686, n1096, n_5249);
  not g10295 (n_5250, n5686);
  and g10296 (n5687, n1100, n_5250);
  not g10297 (n_5251, n5687);
  and g10298 (n5688, n1104, n_5251);
  not g10299 (n_5252, n5688);
  and g10300 (n5689, n1108, n_5252);
  not g10301 (n_5253, n5689);
  and g10302 (n5690, n1112, n_5253);
  not g10303 (n_5254, n5690);
  and g10304 (n5691, n1116, n_5254);
  not g10305 (n_5255, n5691);
  and g10306 (n5692, n1120, n_5255);
  not g10307 (n_5256, n5692);
  and g10308 (n5693, n1124, n_5256);
  not g10309 (n_5257, n5693);
  and g10310 (n5694, n1128, n_5257);
  not g10311 (n_5258, n5694);
  and g10312 (n5695, n1132, n_5258);
  not g10313 (n_5259, n5695);
  and g10314 (n5696, n1136, n_5259);
  not g10315 (n_5260, n5696);
  and g10316 (n5697, n1140, n_5260);
  not g10317 (n_5261, n5697);
  and g10318 (n5698, n1144, n_5261);
  not g10319 (n_5262, n5698);
  and g10320 (n5699, n1148, n_5262);
  not g10321 (n_5263, n5699);
  and g10322 (n5700, n1152, n_5263);
  not g10323 (n_5264, n5700);
  and g10324 (n5701, n1156, n_5264);
  not g10325 (n_5265, n5701);
  and g10326 (n5702, n1160, n_5265);
  not g10327 (n_5266, n5702);
  and g10328 (n5703, n1164, n_5266);
  not g10329 (n_5267, n5703);
  and g10330 (n5704, n1168, n_5267);
  not g10331 (n_5268, n5704);
  and g10332 (n5705, n1172, n_5268);
  not g10333 (n_5269, n5705);
  and g10334 (n5706, n1176, n_5269);
  not g10335 (n_5270, n5706);
  and g10336 (n5707, n1180, n_5270);
  not g10337 (n_5271, n5707);
  and g10338 (n5708, n1184, n_5271);
  not g10339 (n_5272, n5708);
  and g10340 (n5709, n1188, n_5272);
  and g10341 (n5710, \req[52] , n_915);
  not g10342 (n_5273, n5709);
  and g10343 (\grant[52] , n_5273, n5710);
  not g10344 (n_5274, n527);
  and g10345 (n5712, n_5274, n1199);
  not g10346 (n_5275, n5712);
  and g10347 (n5713, n1204, n_5275);
  not g10348 (n_5276, n5713);
  and g10349 (n5714, n1208, n_5276);
  not g10350 (n_5277, n5714);
  and g10351 (n5715, n1212, n_5277);
  not g10352 (n_5278, n5715);
  and g10353 (n5716, n1216, n_5278);
  not g10354 (n_5279, n5716);
  and g10355 (n5717, n1220, n_5279);
  not g10356 (n_5280, n5717);
  and g10357 (n5718, n1224, n_5280);
  not g10358 (n_5281, n5718);
  and g10359 (n5719, n1228, n_5281);
  not g10360 (n_5282, n5719);
  and g10361 (n5720, n1232, n_5282);
  not g10362 (n_5283, n5720);
  and g10363 (n5721, n1236, n_5283);
  not g10364 (n_5284, n5721);
  and g10365 (n5722, n1240, n_5284);
  not g10366 (n_5285, n5722);
  and g10367 (n5723, n1244, n_5285);
  not g10368 (n_5286, n5723);
  and g10369 (n5724, n1248, n_5286);
  not g10370 (n_5287, n5724);
  and g10371 (n5725, n1252, n_5287);
  not g10372 (n_5288, n5725);
  and g10373 (n5726, n1256, n_5288);
  not g10374 (n_5289, n5726);
  and g10375 (n5727, n1260, n_5289);
  not g10376 (n_5290, n5727);
  and g10377 (n5728, n1264, n_5290);
  not g10378 (n_5291, n5728);
  and g10379 (n5729, n1268, n_5291);
  not g10380 (n_5292, n5729);
  and g10381 (n5730, n1272, n_5292);
  not g10382 (n_5293, n5730);
  and g10383 (n5731, n1276, n_5293);
  not g10384 (n_5294, n5731);
  and g10385 (n5732, n1280, n_5294);
  not g10386 (n_5295, n5732);
  and g10387 (n5733, n1284, n_5295);
  not g10388 (n_5296, n5733);
  and g10389 (n5734, n1288, n_5296);
  not g10390 (n_5297, n5734);
  and g10391 (n5735, n1292, n_5297);
  not g10392 (n_5298, n5735);
  and g10393 (n5736, n1296, n_5298);
  not g10394 (n_5299, n5736);
  and g10395 (n5737, n1300, n_5299);
  not g10396 (n_5300, n5737);
  and g10397 (n5738, n1304, n_5300);
  not g10398 (n_5301, n5738);
  and g10399 (n5739, n1308, n_5301);
  not g10400 (n_5302, n5739);
  and g10401 (n5740, n1312, n_5302);
  not g10402 (n_5303, n5740);
  and g10403 (n5741, n1316, n_5303);
  not g10404 (n_5304, n5741);
  and g10405 (n5742, n1320, n_5304);
  not g10406 (n_5305, n5742);
  and g10407 (n5743, n1324, n_5305);
  not g10408 (n_5306, n5743);
  and g10409 (n5744, n1328, n_5306);
  not g10410 (n_5307, n5744);
  and g10411 (n5745, n1332, n_5307);
  not g10412 (n_5308, n5745);
  and g10413 (n5746, n1336, n_5308);
  not g10414 (n_5309, n5746);
  and g10415 (n5747, n1340, n_5309);
  not g10416 (n_5310, n5747);
  and g10417 (n5748, n1344, n_5310);
  not g10418 (n_5311, n5748);
  and g10419 (n5749, n1348, n_5311);
  not g10420 (n_5312, n5749);
  and g10421 (n5750, n1352, n_5312);
  not g10422 (n_5313, n5750);
  and g10423 (n5751, n1356, n_5313);
  not g10424 (n_5314, n5751);
  and g10425 (n5752, n1360, n_5314);
  not g10426 (n_5315, n5752);
  and g10427 (n5753, n1364, n_5315);
  not g10428 (n_5316, n5753);
  and g10429 (n5754, n1368, n_5316);
  not g10430 (n_5317, n5754);
  and g10431 (n5755, n1372, n_5317);
  not g10432 (n_5318, n5755);
  and g10433 (n5756, n1376, n_5318);
  not g10434 (n_5319, n5756);
  and g10435 (n5757, n1380, n_5319);
  not g10436 (n_5320, n5757);
  and g10437 (n5758, n1384, n_5320);
  not g10438 (n_5321, n5758);
  and g10439 (n5759, n1388, n_5321);
  not g10440 (n_5322, n5759);
  and g10441 (n5760, n1392, n_5322);
  not g10442 (n_5323, n5760);
  and g10443 (n5761, n1396, n_5323);
  not g10444 (n_5324, n5761);
  and g10445 (n5762, n1663, n_5324);
  not g10446 (n_5325, n5762);
  and g10447 (n5763, n392, n_5325);
  not g10448 (n_5326, n5763);
  and g10449 (n5764, n396, n_5326);
  not g10450 (n_5327, n5764);
  and g10451 (n5765, n400, n_5327);
  not g10452 (n_5328, n5765);
  and g10453 (n5766, n404, n_5328);
  not g10454 (n_5329, n5766);
  and g10455 (n5767, n408, n_5329);
  not g10456 (n_5330, n5767);
  and g10457 (n5768, n412, n_5330);
  not g10458 (n_5331, n5768);
  and g10459 (n5769, n416, n_5331);
  not g10460 (n_5332, n5769);
  and g10461 (n5770, n420, n_5332);
  not g10462 (n_5333, n5770);
  and g10463 (n5771, n424, n_5333);
  not g10464 (n_5334, n5771);
  and g10465 (n5772, n428, n_5334);
  not g10466 (n_5335, n5772);
  and g10467 (n5773, n432, n_5335);
  not g10468 (n_5336, n5773);
  and g10469 (n5774, n436, n_5336);
  not g10470 (n_5337, n5774);
  and g10471 (n5775, n440, n_5337);
  not g10472 (n_5338, n5775);
  and g10473 (n5776, n444, n_5338);
  not g10474 (n_5339, n5776);
  and g10475 (n5777, n448, n_5339);
  not g10476 (n_5340, n5777);
  and g10477 (n5778, n452, n_5340);
  not g10478 (n_5341, n5778);
  and g10479 (n5779, n456, n_5341);
  not g10480 (n_5342, n5779);
  and g10481 (n5780, n460, n_5342);
  not g10482 (n_5343, n5780);
  and g10483 (n5781, n464, n_5343);
  not g10484 (n_5344, n5781);
  and g10485 (n5782, n468, n_5344);
  not g10486 (n_5345, n5782);
  and g10487 (n5783, n472, n_5345);
  not g10488 (n_5346, n5783);
  and g10489 (n5784, n476, n_5346);
  not g10490 (n_5347, n5784);
  and g10491 (n5785, n480, n_5347);
  not g10492 (n_5348, n5785);
  and g10493 (n5786, n484, n_5348);
  not g10494 (n_5349, n5786);
  and g10495 (n5787, n488, n_5349);
  not g10496 (n_5350, n5787);
  and g10497 (n5788, n492, n_5350);
  not g10498 (n_5351, n5788);
  and g10499 (n5789, n496, n_5351);
  not g10500 (n_5352, n5789);
  and g10501 (n5790, n500, n_5352);
  not g10502 (n_5353, n5790);
  and g10503 (n5791, n504, n_5353);
  not g10504 (n_5354, n5791);
  and g10505 (n5792, n508, n_5354);
  not g10506 (n_5355, n5792);
  and g10507 (n5793, n512, n_5355);
  not g10508 (n_5356, n5793);
  and g10509 (n5794, n516, n_5356);
  not g10510 (n_5357, n5794);
  and g10511 (n5795, n520, n_5357);
  and g10512 (n5796, \req[53] , n_248);
  not g10513 (n_5358, n5795);
  and g10514 (\grant[53] , n_5358, n5796);
  not g10515 (n_5359, n866);
  and g10516 (n5798, n531, n_5359);
  not g10517 (n_5360, n5798);
  and g10518 (n5799, n536, n_5360);
  not g10519 (n_5361, n5799);
  and g10520 (n5800, n540, n_5361);
  not g10521 (n_5362, n5800);
  and g10522 (n5801, n544, n_5362);
  not g10523 (n_5363, n5801);
  and g10524 (n5802, n548, n_5363);
  not g10525 (n_5364, n5802);
  and g10526 (n5803, n552, n_5364);
  not g10527 (n_5365, n5803);
  and g10528 (n5804, n556, n_5365);
  not g10529 (n_5366, n5804);
  and g10530 (n5805, n560, n_5366);
  not g10531 (n_5367, n5805);
  and g10532 (n5806, n564, n_5367);
  not g10533 (n_5368, n5806);
  and g10534 (n5807, n568, n_5368);
  not g10535 (n_5369, n5807);
  and g10536 (n5808, n572, n_5369);
  not g10537 (n_5370, n5808);
  and g10538 (n5809, n576, n_5370);
  not g10539 (n_5371, n5809);
  and g10540 (n5810, n580, n_5371);
  not g10541 (n_5372, n5810);
  and g10542 (n5811, n584, n_5372);
  not g10543 (n_5373, n5811);
  and g10544 (n5812, n588, n_5373);
  not g10545 (n_5374, n5812);
  and g10546 (n5813, n592, n_5374);
  not g10547 (n_5375, n5813);
  and g10548 (n5814, n596, n_5375);
  not g10549 (n_5376, n5814);
  and g10550 (n5815, n600, n_5376);
  not g10551 (n_5377, n5815);
  and g10552 (n5816, n604, n_5377);
  not g10553 (n_5378, n5816);
  and g10554 (n5817, n608, n_5378);
  not g10555 (n_5379, n5817);
  and g10556 (n5818, n612, n_5379);
  not g10557 (n_5380, n5818);
  and g10558 (n5819, n616, n_5380);
  not g10559 (n_5381, n5819);
  and g10560 (n5820, n620, n_5381);
  not g10561 (n_5382, n5820);
  and g10562 (n5821, n624, n_5382);
  not g10563 (n_5383, n5821);
  and g10564 (n5822, n628, n_5383);
  not g10565 (n_5384, n5822);
  and g10566 (n5823, n632, n_5384);
  not g10567 (n_5385, n5823);
  and g10568 (n5824, n636, n_5385);
  not g10569 (n_5386, n5824);
  and g10570 (n5825, n640, n_5386);
  not g10571 (n_5387, n5825);
  and g10572 (n5826, n644, n_5387);
  not g10573 (n_5388, n5826);
  and g10574 (n5827, n648, n_5388);
  not g10575 (n_5389, n5827);
  and g10576 (n5828, n652, n_5389);
  not g10577 (n_5390, n5828);
  and g10578 (n5829, n656, n_5390);
  not g10579 (n_5391, n5829);
  and g10580 (n5830, n660, n_5391);
  not g10581 (n_5392, n5830);
  and g10582 (n5831, n664, n_5392);
  not g10583 (n_5393, n5831);
  and g10584 (n5832, n668, n_5393);
  not g10585 (n_5394, n5832);
  and g10586 (n5833, n672, n_5394);
  not g10587 (n_5395, n5833);
  and g10588 (n5834, n676, n_5395);
  not g10589 (n_5396, n5834);
  and g10590 (n5835, n680, n_5396);
  not g10591 (n_5397, n5835);
  and g10592 (n5836, n684, n_5397);
  not g10593 (n_5398, n5836);
  and g10594 (n5837, n688, n_5398);
  not g10595 (n_5399, n5837);
  and g10596 (n5838, n692, n_5399);
  not g10597 (n_5400, n5838);
  and g10598 (n5839, n696, n_5400);
  not g10599 (n_5401, n5839);
  and g10600 (n5840, n700, n_5401);
  not g10601 (n_5402, n5840);
  and g10602 (n5841, n704, n_5402);
  not g10603 (n_5403, n5841);
  and g10604 (n5842, n708, n_5403);
  not g10605 (n_5404, n5842);
  and g10606 (n5843, n712, n_5404);
  not g10607 (n_5405, n5843);
  and g10608 (n5844, n716, n_5405);
  not g10609 (n_5406, n5844);
  and g10610 (n5845, n720, n_5406);
  not g10611 (n_5407, n5845);
  and g10612 (n5846, n1484, n_5407);
  not g10613 (n_5408, n5846);
  and g10614 (n5847, n1486, n_5408);
  not g10615 (n_5409, n5847);
  and g10616 (n5848, n1750, n_5409);
  not g10617 (n_5410, n5848);
  and g10618 (n5849, n731, n_5410);
  not g10619 (n_5411, n5849);
  and g10620 (n5850, n735, n_5411);
  not g10621 (n_5412, n5850);
  and g10622 (n5851, n739, n_5412);
  not g10623 (n_5413, n5851);
  and g10624 (n5852, n743, n_5413);
  not g10625 (n_5414, n5852);
  and g10626 (n5853, n747, n_5414);
  not g10627 (n_5415, n5853);
  and g10628 (n5854, n751, n_5415);
  not g10629 (n_5416, n5854);
  and g10630 (n5855, n755, n_5416);
  not g10631 (n_5417, n5855);
  and g10632 (n5856, n759, n_5417);
  not g10633 (n_5418, n5856);
  and g10634 (n5857, n763, n_5418);
  not g10635 (n_5419, n5857);
  and g10636 (n5858, n767, n_5419);
  not g10637 (n_5420, n5858);
  and g10638 (n5859, n771, n_5420);
  not g10639 (n_5421, n5859);
  and g10640 (n5860, n775, n_5421);
  not g10641 (n_5422, n5860);
  and g10642 (n5861, n779, n_5422);
  not g10643 (n_5423, n5861);
  and g10644 (n5862, n783, n_5423);
  not g10645 (n_5424, n5862);
  and g10646 (n5863, n787, n_5424);
  not g10647 (n_5425, n5863);
  and g10648 (n5864, n791, n_5425);
  not g10649 (n_5426, n5864);
  and g10650 (n5865, n795, n_5426);
  not g10651 (n_5427, n5865);
  and g10652 (n5866, n799, n_5427);
  not g10653 (n_5428, n5866);
  and g10654 (n5867, n803, n_5428);
  not g10655 (n_5429, n5867);
  and g10656 (n5868, n807, n_5429);
  not g10657 (n_5430, n5868);
  and g10658 (n5869, n811, n_5430);
  not g10659 (n_5431, n5869);
  and g10660 (n5870, n815, n_5431);
  not g10661 (n_5432, n5870);
  and g10662 (n5871, n819, n_5432);
  not g10663 (n_5433, n5871);
  and g10664 (n5872, n823, n_5433);
  not g10665 (n_5434, n5872);
  and g10666 (n5873, n827, n_5434);
  not g10667 (n_5435, n5873);
  and g10668 (n5874, n831, n_5435);
  not g10669 (n_5436, n5874);
  and g10670 (n5875, n835, n_5436);
  not g10671 (n_5437, n5875);
  and g10672 (n5876, n839, n_5437);
  not g10673 (n_5438, n5876);
  and g10674 (n5877, n843, n_5438);
  not g10675 (n_5439, n5877);
  and g10676 (n5878, n847, n_5439);
  not g10677 (n_5440, n5878);
  and g10678 (n5879, n851, n_5440);
  not g10679 (n_5441, n5879);
  and g10680 (n5880, n855, n_5441);
  not g10681 (n_5442, n5880);
  and g10682 (n5881, n859, n_5442);
  and g10683 (n5882, \req[54] , n_701);
  not g10684 (n_5443, n5881);
  and g10685 (\grant[54] , n_5443, n5882);
  not g10686 (n_5444, n1203);
  and g10687 (n5884, n870, n_5444);
  not g10688 (n_5445, n5884);
  and g10689 (n5885, n875, n_5445);
  not g10690 (n_5446, n5885);
  and g10691 (n5886, n879, n_5446);
  not g10692 (n_5447, n5886);
  and g10693 (n5887, n883, n_5447);
  not g10694 (n_5448, n5887);
  and g10695 (n5888, n887, n_5448);
  not g10696 (n_5449, n5888);
  and g10697 (n5889, n891, n_5449);
  not g10698 (n_5450, n5889);
  and g10699 (n5890, n895, n_5450);
  not g10700 (n_5451, n5890);
  and g10701 (n5891, n899, n_5451);
  not g10702 (n_5452, n5891);
  and g10703 (n5892, n903, n_5452);
  not g10704 (n_5453, n5892);
  and g10705 (n5893, n907, n_5453);
  not g10706 (n_5454, n5893);
  and g10707 (n5894, n911, n_5454);
  not g10708 (n_5455, n5894);
  and g10709 (n5895, n915, n_5455);
  not g10710 (n_5456, n5895);
  and g10711 (n5896, n919, n_5456);
  not g10712 (n_5457, n5896);
  and g10713 (n5897, n923, n_5457);
  not g10714 (n_5458, n5897);
  and g10715 (n5898, n927, n_5458);
  not g10716 (n_5459, n5898);
  and g10717 (n5899, n931, n_5459);
  not g10718 (n_5460, n5899);
  and g10719 (n5900, n935, n_5460);
  not g10720 (n_5461, n5900);
  and g10721 (n5901, n939, n_5461);
  not g10722 (n_5462, n5901);
  and g10723 (n5902, n943, n_5462);
  not g10724 (n_5463, n5902);
  and g10725 (n5903, n947, n_5463);
  not g10726 (n_5464, n5903);
  and g10727 (n5904, n951, n_5464);
  not g10728 (n_5465, n5904);
  and g10729 (n5905, n955, n_5465);
  not g10730 (n_5466, n5905);
  and g10731 (n5906, n959, n_5466);
  not g10732 (n_5467, n5906);
  and g10733 (n5907, n963, n_5467);
  not g10734 (n_5468, n5907);
  and g10735 (n5908, n967, n_5468);
  not g10736 (n_5469, n5908);
  and g10737 (n5909, n971, n_5469);
  not g10738 (n_5470, n5909);
  and g10739 (n5910, n975, n_5470);
  not g10740 (n_5471, n5910);
  and g10741 (n5911, n979, n_5471);
  not g10742 (n_5472, n5911);
  and g10743 (n5912, n983, n_5472);
  not g10744 (n_5473, n5912);
  and g10745 (n5913, n987, n_5473);
  not g10746 (n_5474, n5913);
  and g10747 (n5914, n991, n_5474);
  not g10748 (n_5475, n5914);
  and g10749 (n5915, n995, n_5475);
  not g10750 (n_5476, n5915);
  and g10751 (n5916, n999, n_5476);
  not g10752 (n_5477, n5916);
  and g10753 (n5917, n1003, n_5477);
  not g10754 (n_5478, n5917);
  and g10755 (n5918, n1007, n_5478);
  not g10756 (n_5479, n5918);
  and g10757 (n5919, n1011, n_5479);
  not g10758 (n_5480, n5919);
  and g10759 (n5920, n1015, n_5480);
  not g10760 (n_5481, n5920);
  and g10761 (n5921, n1019, n_5481);
  not g10762 (n_5482, n5921);
  and g10763 (n5922, n1023, n_5482);
  not g10764 (n_5483, n5922);
  and g10765 (n5923, n1027, n_5483);
  not g10766 (n_5484, n5923);
  and g10767 (n5924, n1031, n_5484);
  not g10768 (n_5485, n5924);
  and g10769 (n5925, n1035, n_5485);
  not g10770 (n_5486, n5925);
  and g10771 (n5926, n1039, n_5486);
  not g10772 (n_5487, n5926);
  and g10773 (n5927, n1043, n_5487);
  not g10774 (n_5488, n5927);
  and g10775 (n5928, n1047, n_5488);
  not g10776 (n_5489, n5928);
  and g10777 (n5929, n1051, n_5489);
  not g10778 (n_5490, n5929);
  and g10779 (n5930, n1055, n_5490);
  not g10780 (n_5491, n5930);
  and g10781 (n5931, n1059, n_5491);
  not g10782 (n_5492, n5931);
  and g10783 (n5932, n1574, n_5492);
  not g10784 (n_5493, n5932);
  and g10785 (n5933, n1576, n_5493);
  not g10786 (n_5494, n5933);
  and g10787 (n5934, n1837, n_5494);
  not g10788 (n_5495, n5934);
  and g10789 (n5935, n1068, n_5495);
  not g10790 (n_5496, n5935);
  and g10791 (n5936, n1072, n_5496);
  not g10792 (n_5497, n5936);
  and g10793 (n5937, n1076, n_5497);
  not g10794 (n_5498, n5937);
  and g10795 (n5938, n1080, n_5498);
  not g10796 (n_5499, n5938);
  and g10797 (n5939, n1084, n_5499);
  not g10798 (n_5500, n5939);
  and g10799 (n5940, n1088, n_5500);
  not g10800 (n_5501, n5940);
  and g10801 (n5941, n1092, n_5501);
  not g10802 (n_5502, n5941);
  and g10803 (n5942, n1096, n_5502);
  not g10804 (n_5503, n5942);
  and g10805 (n5943, n1100, n_5503);
  not g10806 (n_5504, n5943);
  and g10807 (n5944, n1104, n_5504);
  not g10808 (n_5505, n5944);
  and g10809 (n5945, n1108, n_5505);
  not g10810 (n_5506, n5945);
  and g10811 (n5946, n1112, n_5506);
  not g10812 (n_5507, n5946);
  and g10813 (n5947, n1116, n_5507);
  not g10814 (n_5508, n5947);
  and g10815 (n5948, n1120, n_5508);
  not g10816 (n_5509, n5948);
  and g10817 (n5949, n1124, n_5509);
  not g10818 (n_5510, n5949);
  and g10819 (n5950, n1128, n_5510);
  not g10820 (n_5511, n5950);
  and g10821 (n5951, n1132, n_5511);
  not g10822 (n_5512, n5951);
  and g10823 (n5952, n1136, n_5512);
  not g10824 (n_5513, n5952);
  and g10825 (n5953, n1140, n_5513);
  not g10826 (n_5514, n5953);
  and g10827 (n5954, n1144, n_5514);
  not g10828 (n_5515, n5954);
  and g10829 (n5955, n1148, n_5515);
  not g10830 (n_5516, n5955);
  and g10831 (n5956, n1152, n_5516);
  not g10832 (n_5517, n5956);
  and g10833 (n5957, n1156, n_5517);
  not g10834 (n_5518, n5957);
  and g10835 (n5958, n1160, n_5518);
  not g10836 (n_5519, n5958);
  and g10837 (n5959, n1164, n_5519);
  not g10838 (n_5520, n5959);
  and g10839 (n5960, n1168, n_5520);
  not g10840 (n_5521, n5960);
  and g10841 (n5961, n1172, n_5521);
  not g10842 (n_5522, n5961);
  and g10843 (n5962, n1176, n_5522);
  not g10844 (n_5523, n5962);
  and g10845 (n5963, n1180, n_5523);
  not g10846 (n_5524, n5963);
  and g10847 (n5964, n1184, n_5524);
  not g10848 (n_5525, n5964);
  and g10849 (n5965, n1188, n_5525);
  not g10850 (n_5526, n5965);
  and g10851 (n5966, n1192, n_5526);
  not g10852 (n_5527, n5966);
  and g10853 (n5967, n1196, n_5527);
  and g10854 (n5968, \req[55] , n_919);
  not g10855 (n_5528, n5967);
  and g10856 (\grant[55] , n_5528, n5968);
  not g10857 (n_5529, n535);
  and g10858 (n5970, n_5529, n1207);
  not g10859 (n_5530, n5970);
  and g10860 (n5971, n1212, n_5530);
  not g10861 (n_5531, n5971);
  and g10862 (n5972, n1216, n_5531);
  not g10863 (n_5532, n5972);
  and g10864 (n5973, n1220, n_5532);
  not g10865 (n_5533, n5973);
  and g10866 (n5974, n1224, n_5533);
  not g10867 (n_5534, n5974);
  and g10868 (n5975, n1228, n_5534);
  not g10869 (n_5535, n5975);
  and g10870 (n5976, n1232, n_5535);
  not g10871 (n_5536, n5976);
  and g10872 (n5977, n1236, n_5536);
  not g10873 (n_5537, n5977);
  and g10874 (n5978, n1240, n_5537);
  not g10875 (n_5538, n5978);
  and g10876 (n5979, n1244, n_5538);
  not g10877 (n_5539, n5979);
  and g10878 (n5980, n1248, n_5539);
  not g10879 (n_5540, n5980);
  and g10880 (n5981, n1252, n_5540);
  not g10881 (n_5541, n5981);
  and g10882 (n5982, n1256, n_5541);
  not g10883 (n_5542, n5982);
  and g10884 (n5983, n1260, n_5542);
  not g10885 (n_5543, n5983);
  and g10886 (n5984, n1264, n_5543);
  not g10887 (n_5544, n5984);
  and g10888 (n5985, n1268, n_5544);
  not g10889 (n_5545, n5985);
  and g10890 (n5986, n1272, n_5545);
  not g10891 (n_5546, n5986);
  and g10892 (n5987, n1276, n_5546);
  not g10893 (n_5547, n5987);
  and g10894 (n5988, n1280, n_5547);
  not g10895 (n_5548, n5988);
  and g10896 (n5989, n1284, n_5548);
  not g10897 (n_5549, n5989);
  and g10898 (n5990, n1288, n_5549);
  not g10899 (n_5550, n5990);
  and g10900 (n5991, n1292, n_5550);
  not g10901 (n_5551, n5991);
  and g10902 (n5992, n1296, n_5551);
  not g10903 (n_5552, n5992);
  and g10904 (n5993, n1300, n_5552);
  not g10905 (n_5553, n5993);
  and g10906 (n5994, n1304, n_5553);
  not g10907 (n_5554, n5994);
  and g10908 (n5995, n1308, n_5554);
  not g10909 (n_5555, n5995);
  and g10910 (n5996, n1312, n_5555);
  not g10911 (n_5556, n5996);
  and g10912 (n5997, n1316, n_5556);
  not g10913 (n_5557, n5997);
  and g10914 (n5998, n1320, n_5557);
  not g10915 (n_5558, n5998);
  and g10916 (n5999, n1324, n_5558);
  not g10917 (n_5559, n5999);
  and g10918 (n6000, n1328, n_5559);
  not g10919 (n_5560, n6000);
  and g10920 (n6001, n1332, n_5560);
  not g10921 (n_5561, n6001);
  and g10922 (n6002, n1336, n_5561);
  not g10923 (n_5562, n6002);
  and g10924 (n6003, n1340, n_5562);
  not g10925 (n_5563, n6003);
  and g10926 (n6004, n1344, n_5563);
  not g10927 (n_5564, n6004);
  and g10928 (n6005, n1348, n_5564);
  not g10929 (n_5565, n6005);
  and g10930 (n6006, n1352, n_5565);
  not g10931 (n_5566, n6006);
  and g10932 (n6007, n1356, n_5566);
  not g10933 (n_5567, n6007);
  and g10934 (n6008, n1360, n_5567);
  not g10935 (n_5568, n6008);
  and g10936 (n6009, n1364, n_5568);
  not g10937 (n_5569, n6009);
  and g10938 (n6010, n1368, n_5569);
  not g10939 (n_5570, n6010);
  and g10940 (n6011, n1372, n_5570);
  not g10941 (n_5571, n6011);
  and g10942 (n6012, n1376, n_5571);
  not g10943 (n_5572, n6012);
  and g10944 (n6013, n1380, n_5572);
  not g10945 (n_5573, n6013);
  and g10946 (n6014, n1384, n_5573);
  not g10947 (n_5574, n6014);
  and g10948 (n6015, n1388, n_5574);
  not g10949 (n_5575, n6015);
  and g10950 (n6016, n1392, n_5575);
  not g10951 (n_5576, n6016);
  and g10952 (n6017, n1396, n_5576);
  not g10953 (n_5577, n6017);
  and g10954 (n6018, n1663, n_5577);
  not g10955 (n_5578, n6018);
  and g10956 (n6019, n392, n_5578);
  not g10957 (n_5579, n6019);
  and g10958 (n6020, n396, n_5579);
  not g10959 (n_5580, n6020);
  and g10960 (n6021, n400, n_5580);
  not g10961 (n_5581, n6021);
  and g10962 (n6022, n404, n_5581);
  not g10963 (n_5582, n6022);
  and g10964 (n6023, n408, n_5582);
  not g10965 (n_5583, n6023);
  and g10966 (n6024, n412, n_5583);
  not g10967 (n_5584, n6024);
  and g10968 (n6025, n416, n_5584);
  not g10969 (n_5585, n6025);
  and g10970 (n6026, n420, n_5585);
  not g10971 (n_5586, n6026);
  and g10972 (n6027, n424, n_5586);
  not g10973 (n_5587, n6027);
  and g10974 (n6028, n428, n_5587);
  not g10975 (n_5588, n6028);
  and g10976 (n6029, n432, n_5588);
  not g10977 (n_5589, n6029);
  and g10978 (n6030, n436, n_5589);
  not g10979 (n_5590, n6030);
  and g10980 (n6031, n440, n_5590);
  not g10981 (n_5591, n6031);
  and g10982 (n6032, n444, n_5591);
  not g10983 (n_5592, n6032);
  and g10984 (n6033, n448, n_5592);
  not g10985 (n_5593, n6033);
  and g10986 (n6034, n452, n_5593);
  not g10987 (n_5594, n6034);
  and g10988 (n6035, n456, n_5594);
  not g10989 (n_5595, n6035);
  and g10990 (n6036, n460, n_5595);
  not g10991 (n_5596, n6036);
  and g10992 (n6037, n464, n_5596);
  not g10993 (n_5597, n6037);
  and g10994 (n6038, n468, n_5597);
  not g10995 (n_5598, n6038);
  and g10996 (n6039, n472, n_5598);
  not g10997 (n_5599, n6039);
  and g10998 (n6040, n476, n_5599);
  not g10999 (n_5600, n6040);
  and g11000 (n6041, n480, n_5600);
  not g11001 (n_5601, n6041);
  and g11002 (n6042, n484, n_5601);
  not g11003 (n_5602, n6042);
  and g11004 (n6043, n488, n_5602);
  not g11005 (n_5603, n6043);
  and g11006 (n6044, n492, n_5603);
  not g11007 (n_5604, n6044);
  and g11008 (n6045, n496, n_5604);
  not g11009 (n_5605, n6045);
  and g11010 (n6046, n500, n_5605);
  not g11011 (n_5606, n6046);
  and g11012 (n6047, n504, n_5606);
  not g11013 (n_5607, n6047);
  and g11014 (n6048, n508, n_5607);
  not g11015 (n_5608, n6048);
  and g11016 (n6049, n512, n_5608);
  not g11017 (n_5609, n6049);
  and g11018 (n6050, n516, n_5609);
  not g11019 (n_5610, n6050);
  and g11020 (n6051, n520, n_5610);
  not g11021 (n_5611, n6051);
  and g11022 (n6052, n524, n_5611);
  not g11023 (n_5612, n6052);
  and g11024 (n6053, n528, n_5612);
  and g11025 (n6054, \req[56] , n_262);
  not g11026 (n_5613, n6053);
  and g11027 (\grant[56] , n_5613, n6054);
  not g11028 (n_5614, n874);
  and g11029 (n6056, n539, n_5614);
  not g11030 (n_5615, n6056);
  and g11031 (n6057, n544, n_5615);
  not g11032 (n_5616, n6057);
  and g11033 (n6058, n548, n_5616);
  not g11034 (n_5617, n6058);
  and g11035 (n6059, n552, n_5617);
  not g11036 (n_5618, n6059);
  and g11037 (n6060, n556, n_5618);
  not g11038 (n_5619, n6060);
  and g11039 (n6061, n560, n_5619);
  not g11040 (n_5620, n6061);
  and g11041 (n6062, n564, n_5620);
  not g11042 (n_5621, n6062);
  and g11043 (n6063, n568, n_5621);
  not g11044 (n_5622, n6063);
  and g11045 (n6064, n572, n_5622);
  not g11046 (n_5623, n6064);
  and g11047 (n6065, n576, n_5623);
  not g11048 (n_5624, n6065);
  and g11049 (n6066, n580, n_5624);
  not g11050 (n_5625, n6066);
  and g11051 (n6067, n584, n_5625);
  not g11052 (n_5626, n6067);
  and g11053 (n6068, n588, n_5626);
  not g11054 (n_5627, n6068);
  and g11055 (n6069, n592, n_5627);
  not g11056 (n_5628, n6069);
  and g11057 (n6070, n596, n_5628);
  not g11058 (n_5629, n6070);
  and g11059 (n6071, n600, n_5629);
  not g11060 (n_5630, n6071);
  and g11061 (n6072, n604, n_5630);
  not g11062 (n_5631, n6072);
  and g11063 (n6073, n608, n_5631);
  not g11064 (n_5632, n6073);
  and g11065 (n6074, n612, n_5632);
  not g11066 (n_5633, n6074);
  and g11067 (n6075, n616, n_5633);
  not g11068 (n_5634, n6075);
  and g11069 (n6076, n620, n_5634);
  not g11070 (n_5635, n6076);
  and g11071 (n6077, n624, n_5635);
  not g11072 (n_5636, n6077);
  and g11073 (n6078, n628, n_5636);
  not g11074 (n_5637, n6078);
  and g11075 (n6079, n632, n_5637);
  not g11076 (n_5638, n6079);
  and g11077 (n6080, n636, n_5638);
  not g11078 (n_5639, n6080);
  and g11079 (n6081, n640, n_5639);
  not g11080 (n_5640, n6081);
  and g11081 (n6082, n644, n_5640);
  not g11082 (n_5641, n6082);
  and g11083 (n6083, n648, n_5641);
  not g11084 (n_5642, n6083);
  and g11085 (n6084, n652, n_5642);
  not g11086 (n_5643, n6084);
  and g11087 (n6085, n656, n_5643);
  not g11088 (n_5644, n6085);
  and g11089 (n6086, n660, n_5644);
  not g11090 (n_5645, n6086);
  and g11091 (n6087, n664, n_5645);
  not g11092 (n_5646, n6087);
  and g11093 (n6088, n668, n_5646);
  not g11094 (n_5647, n6088);
  and g11095 (n6089, n672, n_5647);
  not g11096 (n_5648, n6089);
  and g11097 (n6090, n676, n_5648);
  not g11098 (n_5649, n6090);
  and g11099 (n6091, n680, n_5649);
  not g11100 (n_5650, n6091);
  and g11101 (n6092, n684, n_5650);
  not g11102 (n_5651, n6092);
  and g11103 (n6093, n688, n_5651);
  not g11104 (n_5652, n6093);
  and g11105 (n6094, n692, n_5652);
  not g11106 (n_5653, n6094);
  and g11107 (n6095, n696, n_5653);
  not g11108 (n_5654, n6095);
  and g11109 (n6096, n700, n_5654);
  not g11110 (n_5655, n6096);
  and g11111 (n6097, n704, n_5655);
  not g11112 (n_5656, n6097);
  and g11113 (n6098, n708, n_5656);
  not g11114 (n_5657, n6098);
  and g11115 (n6099, n712, n_5657);
  not g11116 (n_5658, n6099);
  and g11117 (n6100, n716, n_5658);
  not g11118 (n_5659, n6100);
  and g11119 (n6101, n720, n_5659);
  not g11120 (n_5660, n6101);
  and g11121 (n6102, n1484, n_5660);
  not g11122 (n_5661, n6102);
  and g11123 (n6103, n1486, n_5661);
  not g11124 (n_5662, n6103);
  and g11125 (n6104, n1750, n_5662);
  not g11126 (n_5663, n6104);
  and g11127 (n6105, n731, n_5663);
  not g11128 (n_5664, n6105);
  and g11129 (n6106, n735, n_5664);
  not g11130 (n_5665, n6106);
  and g11131 (n6107, n739, n_5665);
  not g11132 (n_5666, n6107);
  and g11133 (n6108, n743, n_5666);
  not g11134 (n_5667, n6108);
  and g11135 (n6109, n747, n_5667);
  not g11136 (n_5668, n6109);
  and g11137 (n6110, n751, n_5668);
  not g11138 (n_5669, n6110);
  and g11139 (n6111, n755, n_5669);
  not g11140 (n_5670, n6111);
  and g11141 (n6112, n759, n_5670);
  not g11142 (n_5671, n6112);
  and g11143 (n6113, n763, n_5671);
  not g11144 (n_5672, n6113);
  and g11145 (n6114, n767, n_5672);
  not g11146 (n_5673, n6114);
  and g11147 (n6115, n771, n_5673);
  not g11148 (n_5674, n6115);
  and g11149 (n6116, n775, n_5674);
  not g11150 (n_5675, n6116);
  and g11151 (n6117, n779, n_5675);
  not g11152 (n_5676, n6117);
  and g11153 (n6118, n783, n_5676);
  not g11154 (n_5677, n6118);
  and g11155 (n6119, n787, n_5677);
  not g11156 (n_5678, n6119);
  and g11157 (n6120, n791, n_5678);
  not g11158 (n_5679, n6120);
  and g11159 (n6121, n795, n_5679);
  not g11160 (n_5680, n6121);
  and g11161 (n6122, n799, n_5680);
  not g11162 (n_5681, n6122);
  and g11163 (n6123, n803, n_5681);
  not g11164 (n_5682, n6123);
  and g11165 (n6124, n807, n_5682);
  not g11166 (n_5683, n6124);
  and g11167 (n6125, n811, n_5683);
  not g11168 (n_5684, n6125);
  and g11169 (n6126, n815, n_5684);
  not g11170 (n_5685, n6126);
  and g11171 (n6127, n819, n_5685);
  not g11172 (n_5686, n6127);
  and g11173 (n6128, n823, n_5686);
  not g11174 (n_5687, n6128);
  and g11175 (n6129, n827, n_5687);
  not g11176 (n_5688, n6129);
  and g11177 (n6130, n831, n_5688);
  not g11178 (n_5689, n6130);
  and g11179 (n6131, n835, n_5689);
  not g11180 (n_5690, n6131);
  and g11181 (n6132, n839, n_5690);
  not g11182 (n_5691, n6132);
  and g11183 (n6133, n843, n_5691);
  not g11184 (n_5692, n6133);
  and g11185 (n6134, n847, n_5692);
  not g11186 (n_5693, n6134);
  and g11187 (n6135, n851, n_5693);
  not g11188 (n_5694, n6135);
  and g11189 (n6136, n855, n_5694);
  not g11190 (n_5695, n6136);
  and g11191 (n6137, n859, n_5695);
  not g11192 (n_5696, n6137);
  and g11193 (n6138, n863, n_5696);
  not g11194 (n_5697, n6138);
  and g11195 (n6139, n867, n_5697);
  and g11196 (n6140, \req[57] , n_707);
  not g11197 (n_5698, n6139);
  and g11198 (\grant[57] , n_5698, n6140);
  not g11199 (n_5699, n1211);
  and g11200 (n6142, n878, n_5699);
  not g11201 (n_5700, n6142);
  and g11202 (n6143, n883, n_5700);
  not g11203 (n_5701, n6143);
  and g11204 (n6144, n887, n_5701);
  not g11205 (n_5702, n6144);
  and g11206 (n6145, n891, n_5702);
  not g11207 (n_5703, n6145);
  and g11208 (n6146, n895, n_5703);
  not g11209 (n_5704, n6146);
  and g11210 (n6147, n899, n_5704);
  not g11211 (n_5705, n6147);
  and g11212 (n6148, n903, n_5705);
  not g11213 (n_5706, n6148);
  and g11214 (n6149, n907, n_5706);
  not g11215 (n_5707, n6149);
  and g11216 (n6150, n911, n_5707);
  not g11217 (n_5708, n6150);
  and g11218 (n6151, n915, n_5708);
  not g11219 (n_5709, n6151);
  and g11220 (n6152, n919, n_5709);
  not g11221 (n_5710, n6152);
  and g11222 (n6153, n923, n_5710);
  not g11223 (n_5711, n6153);
  and g11224 (n6154, n927, n_5711);
  not g11225 (n_5712, n6154);
  and g11226 (n6155, n931, n_5712);
  not g11227 (n_5713, n6155);
  and g11228 (n6156, n935, n_5713);
  not g11229 (n_5714, n6156);
  and g11230 (n6157, n939, n_5714);
  not g11231 (n_5715, n6157);
  and g11232 (n6158, n943, n_5715);
  not g11233 (n_5716, n6158);
  and g11234 (n6159, n947, n_5716);
  not g11235 (n_5717, n6159);
  and g11236 (n6160, n951, n_5717);
  not g11237 (n_5718, n6160);
  and g11238 (n6161, n955, n_5718);
  not g11239 (n_5719, n6161);
  and g11240 (n6162, n959, n_5719);
  not g11241 (n_5720, n6162);
  and g11242 (n6163, n963, n_5720);
  not g11243 (n_5721, n6163);
  and g11244 (n6164, n967, n_5721);
  not g11245 (n_5722, n6164);
  and g11246 (n6165, n971, n_5722);
  not g11247 (n_5723, n6165);
  and g11248 (n6166, n975, n_5723);
  not g11249 (n_5724, n6166);
  and g11250 (n6167, n979, n_5724);
  not g11251 (n_5725, n6167);
  and g11252 (n6168, n983, n_5725);
  not g11253 (n_5726, n6168);
  and g11254 (n6169, n987, n_5726);
  not g11255 (n_5727, n6169);
  and g11256 (n6170, n991, n_5727);
  not g11257 (n_5728, n6170);
  and g11258 (n6171, n995, n_5728);
  not g11259 (n_5729, n6171);
  and g11260 (n6172, n999, n_5729);
  not g11261 (n_5730, n6172);
  and g11262 (n6173, n1003, n_5730);
  not g11263 (n_5731, n6173);
  and g11264 (n6174, n1007, n_5731);
  not g11265 (n_5732, n6174);
  and g11266 (n6175, n1011, n_5732);
  not g11267 (n_5733, n6175);
  and g11268 (n6176, n1015, n_5733);
  not g11269 (n_5734, n6176);
  and g11270 (n6177, n1019, n_5734);
  not g11271 (n_5735, n6177);
  and g11272 (n6178, n1023, n_5735);
  not g11273 (n_5736, n6178);
  and g11274 (n6179, n1027, n_5736);
  not g11275 (n_5737, n6179);
  and g11276 (n6180, n1031, n_5737);
  not g11277 (n_5738, n6180);
  and g11278 (n6181, n1035, n_5738);
  not g11279 (n_5739, n6181);
  and g11280 (n6182, n1039, n_5739);
  not g11281 (n_5740, n6182);
  and g11282 (n6183, n1043, n_5740);
  not g11283 (n_5741, n6183);
  and g11284 (n6184, n1047, n_5741);
  not g11285 (n_5742, n6184);
  and g11286 (n6185, n1051, n_5742);
  not g11287 (n_5743, n6185);
  and g11288 (n6186, n1055, n_5743);
  not g11289 (n_5744, n6186);
  and g11290 (n6187, n1059, n_5744);
  not g11291 (n_5745, n6187);
  and g11292 (n6188, n1574, n_5745);
  not g11293 (n_5746, n6188);
  and g11294 (n6189, n1576, n_5746);
  not g11295 (n_5747, n6189);
  and g11296 (n6190, n1837, n_5747);
  not g11297 (n_5748, n6190);
  and g11298 (n6191, n1068, n_5748);
  not g11299 (n_5749, n6191);
  and g11300 (n6192, n1072, n_5749);
  not g11301 (n_5750, n6192);
  and g11302 (n6193, n1076, n_5750);
  not g11303 (n_5751, n6193);
  and g11304 (n6194, n1080, n_5751);
  not g11305 (n_5752, n6194);
  and g11306 (n6195, n1084, n_5752);
  not g11307 (n_5753, n6195);
  and g11308 (n6196, n1088, n_5753);
  not g11309 (n_5754, n6196);
  and g11310 (n6197, n1092, n_5754);
  not g11311 (n_5755, n6197);
  and g11312 (n6198, n1096, n_5755);
  not g11313 (n_5756, n6198);
  and g11314 (n6199, n1100, n_5756);
  not g11315 (n_5757, n6199);
  and g11316 (n6200, n1104, n_5757);
  not g11317 (n_5758, n6200);
  and g11318 (n6201, n1108, n_5758);
  not g11319 (n_5759, n6201);
  and g11320 (n6202, n1112, n_5759);
  not g11321 (n_5760, n6202);
  and g11322 (n6203, n1116, n_5760);
  not g11323 (n_5761, n6203);
  and g11324 (n6204, n1120, n_5761);
  not g11325 (n_5762, n6204);
  and g11326 (n6205, n1124, n_5762);
  not g11327 (n_5763, n6205);
  and g11328 (n6206, n1128, n_5763);
  not g11329 (n_5764, n6206);
  and g11330 (n6207, n1132, n_5764);
  not g11331 (n_5765, n6207);
  and g11332 (n6208, n1136, n_5765);
  not g11333 (n_5766, n6208);
  and g11334 (n6209, n1140, n_5766);
  not g11335 (n_5767, n6209);
  and g11336 (n6210, n1144, n_5767);
  not g11337 (n_5768, n6210);
  and g11338 (n6211, n1148, n_5768);
  not g11339 (n_5769, n6211);
  and g11340 (n6212, n1152, n_5769);
  not g11341 (n_5770, n6212);
  and g11342 (n6213, n1156, n_5770);
  not g11343 (n_5771, n6213);
  and g11344 (n6214, n1160, n_5771);
  not g11345 (n_5772, n6214);
  and g11346 (n6215, n1164, n_5772);
  not g11347 (n_5773, n6215);
  and g11348 (n6216, n1168, n_5773);
  not g11349 (n_5774, n6216);
  and g11350 (n6217, n1172, n_5774);
  not g11351 (n_5775, n6217);
  and g11352 (n6218, n1176, n_5775);
  not g11353 (n_5776, n6218);
  and g11354 (n6219, n1180, n_5776);
  not g11355 (n_5777, n6219);
  and g11356 (n6220, n1184, n_5777);
  not g11357 (n_5778, n6220);
  and g11358 (n6221, n1188, n_5778);
  not g11359 (n_5779, n6221);
  and g11360 (n6222, n1192, n_5779);
  not g11361 (n_5780, n6222);
  and g11362 (n6223, n1196, n_5780);
  not g11363 (n_5781, n6223);
  and g11364 (n6224, n1200, n_5781);
  not g11365 (n_5782, n6224);
  and g11366 (n6225, n1204, n_5782);
  and g11367 (n6226, \req[58] , n_923);
  not g11368 (n_5783, n6225);
  and g11369 (\grant[58] , n_5783, n6226);
  not g11370 (n_5784, n543);
  and g11371 (n6228, n_5784, n1215);
  not g11372 (n_5785, n6228);
  and g11373 (n6229, n1220, n_5785);
  not g11374 (n_5786, n6229);
  and g11375 (n6230, n1224, n_5786);
  not g11376 (n_5787, n6230);
  and g11377 (n6231, n1228, n_5787);
  not g11378 (n_5788, n6231);
  and g11379 (n6232, n1232, n_5788);
  not g11380 (n_5789, n6232);
  and g11381 (n6233, n1236, n_5789);
  not g11382 (n_5790, n6233);
  and g11383 (n6234, n1240, n_5790);
  not g11384 (n_5791, n6234);
  and g11385 (n6235, n1244, n_5791);
  not g11386 (n_5792, n6235);
  and g11387 (n6236, n1248, n_5792);
  not g11388 (n_5793, n6236);
  and g11389 (n6237, n1252, n_5793);
  not g11390 (n_5794, n6237);
  and g11391 (n6238, n1256, n_5794);
  not g11392 (n_5795, n6238);
  and g11393 (n6239, n1260, n_5795);
  not g11394 (n_5796, n6239);
  and g11395 (n6240, n1264, n_5796);
  not g11396 (n_5797, n6240);
  and g11397 (n6241, n1268, n_5797);
  not g11398 (n_5798, n6241);
  and g11399 (n6242, n1272, n_5798);
  not g11400 (n_5799, n6242);
  and g11401 (n6243, n1276, n_5799);
  not g11402 (n_5800, n6243);
  and g11403 (n6244, n1280, n_5800);
  not g11404 (n_5801, n6244);
  and g11405 (n6245, n1284, n_5801);
  not g11406 (n_5802, n6245);
  and g11407 (n6246, n1288, n_5802);
  not g11408 (n_5803, n6246);
  and g11409 (n6247, n1292, n_5803);
  not g11410 (n_5804, n6247);
  and g11411 (n6248, n1296, n_5804);
  not g11412 (n_5805, n6248);
  and g11413 (n6249, n1300, n_5805);
  not g11414 (n_5806, n6249);
  and g11415 (n6250, n1304, n_5806);
  not g11416 (n_5807, n6250);
  and g11417 (n6251, n1308, n_5807);
  not g11418 (n_5808, n6251);
  and g11419 (n6252, n1312, n_5808);
  not g11420 (n_5809, n6252);
  and g11421 (n6253, n1316, n_5809);
  not g11422 (n_5810, n6253);
  and g11423 (n6254, n1320, n_5810);
  not g11424 (n_5811, n6254);
  and g11425 (n6255, n1324, n_5811);
  not g11426 (n_5812, n6255);
  and g11427 (n6256, n1328, n_5812);
  not g11428 (n_5813, n6256);
  and g11429 (n6257, n1332, n_5813);
  not g11430 (n_5814, n6257);
  and g11431 (n6258, n1336, n_5814);
  not g11432 (n_5815, n6258);
  and g11433 (n6259, n1340, n_5815);
  not g11434 (n_5816, n6259);
  and g11435 (n6260, n1344, n_5816);
  not g11436 (n_5817, n6260);
  and g11437 (n6261, n1348, n_5817);
  not g11438 (n_5818, n6261);
  and g11439 (n6262, n1352, n_5818);
  not g11440 (n_5819, n6262);
  and g11441 (n6263, n1356, n_5819);
  not g11442 (n_5820, n6263);
  and g11443 (n6264, n1360, n_5820);
  not g11444 (n_5821, n6264);
  and g11445 (n6265, n1364, n_5821);
  not g11446 (n_5822, n6265);
  and g11447 (n6266, n1368, n_5822);
  not g11448 (n_5823, n6266);
  and g11449 (n6267, n1372, n_5823);
  not g11450 (n_5824, n6267);
  and g11451 (n6268, n1376, n_5824);
  not g11452 (n_5825, n6268);
  and g11453 (n6269, n1380, n_5825);
  not g11454 (n_5826, n6269);
  and g11455 (n6270, n1384, n_5826);
  not g11456 (n_5827, n6270);
  and g11457 (n6271, n1388, n_5827);
  not g11458 (n_5828, n6271);
  and g11459 (n6272, n1392, n_5828);
  not g11460 (n_5829, n6272);
  and g11461 (n6273, n1396, n_5829);
  not g11462 (n_5830, n6273);
  and g11463 (n6274, n1663, n_5830);
  not g11464 (n_5831, n6274);
  and g11465 (n6275, n392, n_5831);
  not g11466 (n_5832, n6275);
  and g11467 (n6276, n396, n_5832);
  not g11468 (n_5833, n6276);
  and g11469 (n6277, n400, n_5833);
  not g11470 (n_5834, n6277);
  and g11471 (n6278, n404, n_5834);
  not g11472 (n_5835, n6278);
  and g11473 (n6279, n408, n_5835);
  not g11474 (n_5836, n6279);
  and g11475 (n6280, n412, n_5836);
  not g11476 (n_5837, n6280);
  and g11477 (n6281, n416, n_5837);
  not g11478 (n_5838, n6281);
  and g11479 (n6282, n420, n_5838);
  not g11480 (n_5839, n6282);
  and g11481 (n6283, n424, n_5839);
  not g11482 (n_5840, n6283);
  and g11483 (n6284, n428, n_5840);
  not g11484 (n_5841, n6284);
  and g11485 (n6285, n432, n_5841);
  not g11486 (n_5842, n6285);
  and g11487 (n6286, n436, n_5842);
  not g11488 (n_5843, n6286);
  and g11489 (n6287, n440, n_5843);
  not g11490 (n_5844, n6287);
  and g11491 (n6288, n444, n_5844);
  not g11492 (n_5845, n6288);
  and g11493 (n6289, n448, n_5845);
  not g11494 (n_5846, n6289);
  and g11495 (n6290, n452, n_5846);
  not g11496 (n_5847, n6290);
  and g11497 (n6291, n456, n_5847);
  not g11498 (n_5848, n6291);
  and g11499 (n6292, n460, n_5848);
  not g11500 (n_5849, n6292);
  and g11501 (n6293, n464, n_5849);
  not g11502 (n_5850, n6293);
  and g11503 (n6294, n468, n_5850);
  not g11504 (n_5851, n6294);
  and g11505 (n6295, n472, n_5851);
  not g11506 (n_5852, n6295);
  and g11507 (n6296, n476, n_5852);
  not g11508 (n_5853, n6296);
  and g11509 (n6297, n480, n_5853);
  not g11510 (n_5854, n6297);
  and g11511 (n6298, n484, n_5854);
  not g11512 (n_5855, n6298);
  and g11513 (n6299, n488, n_5855);
  not g11514 (n_5856, n6299);
  and g11515 (n6300, n492, n_5856);
  not g11516 (n_5857, n6300);
  and g11517 (n6301, n496, n_5857);
  not g11518 (n_5858, n6301);
  and g11519 (n6302, n500, n_5858);
  not g11520 (n_5859, n6302);
  and g11521 (n6303, n504, n_5859);
  not g11522 (n_5860, n6303);
  and g11523 (n6304, n508, n_5860);
  not g11524 (n_5861, n6304);
  and g11525 (n6305, n512, n_5861);
  not g11526 (n_5862, n6305);
  and g11527 (n6306, n516, n_5862);
  not g11528 (n_5863, n6306);
  and g11529 (n6307, n520, n_5863);
  not g11530 (n_5864, n6307);
  and g11531 (n6308, n524, n_5864);
  not g11532 (n_5865, n6308);
  and g11533 (n6309, n528, n_5865);
  not g11534 (n_5866, n6309);
  and g11535 (n6310, n532, n_5866);
  not g11536 (n_5867, n6310);
  and g11537 (n6311, n536, n_5867);
  and g11538 (n6312, \req[59] , n_276);
  not g11539 (n_5868, n6311);
  and g11540 (\grant[59] , n_5868, n6312);
  not g11541 (n_5869, n882);
  and g11542 (n6314, n547, n_5869);
  not g11543 (n_5870, n6314);
  and g11544 (n6315, n552, n_5870);
  not g11545 (n_5871, n6315);
  and g11546 (n6316, n556, n_5871);
  not g11547 (n_5872, n6316);
  and g11548 (n6317, n560, n_5872);
  not g11549 (n_5873, n6317);
  and g11550 (n6318, n564, n_5873);
  not g11551 (n_5874, n6318);
  and g11552 (n6319, n568, n_5874);
  not g11553 (n_5875, n6319);
  and g11554 (n6320, n572, n_5875);
  not g11555 (n_5876, n6320);
  and g11556 (n6321, n576, n_5876);
  not g11557 (n_5877, n6321);
  and g11558 (n6322, n580, n_5877);
  not g11559 (n_5878, n6322);
  and g11560 (n6323, n584, n_5878);
  not g11561 (n_5879, n6323);
  and g11562 (n6324, n588, n_5879);
  not g11563 (n_5880, n6324);
  and g11564 (n6325, n592, n_5880);
  not g11565 (n_5881, n6325);
  and g11566 (n6326, n596, n_5881);
  not g11567 (n_5882, n6326);
  and g11568 (n6327, n600, n_5882);
  not g11569 (n_5883, n6327);
  and g11570 (n6328, n604, n_5883);
  not g11571 (n_5884, n6328);
  and g11572 (n6329, n608, n_5884);
  not g11573 (n_5885, n6329);
  and g11574 (n6330, n612, n_5885);
  not g11575 (n_5886, n6330);
  and g11576 (n6331, n616, n_5886);
  not g11577 (n_5887, n6331);
  and g11578 (n6332, n620, n_5887);
  not g11579 (n_5888, n6332);
  and g11580 (n6333, n624, n_5888);
  not g11581 (n_5889, n6333);
  and g11582 (n6334, n628, n_5889);
  not g11583 (n_5890, n6334);
  and g11584 (n6335, n632, n_5890);
  not g11585 (n_5891, n6335);
  and g11586 (n6336, n636, n_5891);
  not g11587 (n_5892, n6336);
  and g11588 (n6337, n640, n_5892);
  not g11589 (n_5893, n6337);
  and g11590 (n6338, n644, n_5893);
  not g11591 (n_5894, n6338);
  and g11592 (n6339, n648, n_5894);
  not g11593 (n_5895, n6339);
  and g11594 (n6340, n652, n_5895);
  not g11595 (n_5896, n6340);
  and g11596 (n6341, n656, n_5896);
  not g11597 (n_5897, n6341);
  and g11598 (n6342, n660, n_5897);
  not g11599 (n_5898, n6342);
  and g11600 (n6343, n664, n_5898);
  not g11601 (n_5899, n6343);
  and g11602 (n6344, n668, n_5899);
  not g11603 (n_5900, n6344);
  and g11604 (n6345, n672, n_5900);
  not g11605 (n_5901, n6345);
  and g11606 (n6346, n676, n_5901);
  not g11607 (n_5902, n6346);
  and g11608 (n6347, n680, n_5902);
  not g11609 (n_5903, n6347);
  and g11610 (n6348, n684, n_5903);
  not g11611 (n_5904, n6348);
  and g11612 (n6349, n688, n_5904);
  not g11613 (n_5905, n6349);
  and g11614 (n6350, n692, n_5905);
  not g11615 (n_5906, n6350);
  and g11616 (n6351, n696, n_5906);
  not g11617 (n_5907, n6351);
  and g11618 (n6352, n700, n_5907);
  not g11619 (n_5908, n6352);
  and g11620 (n6353, n704, n_5908);
  not g11621 (n_5909, n6353);
  and g11622 (n6354, n708, n_5909);
  not g11623 (n_5910, n6354);
  and g11624 (n6355, n712, n_5910);
  not g11625 (n_5911, n6355);
  and g11626 (n6356, n716, n_5911);
  not g11627 (n_5912, n6356);
  and g11628 (n6357, n720, n_5912);
  not g11629 (n_5913, n6357);
  and g11630 (n6358, n1484, n_5913);
  not g11631 (n_5914, n6358);
  and g11632 (n6359, n1486, n_5914);
  not g11633 (n_5915, n6359);
  and g11634 (n6360, n1750, n_5915);
  not g11635 (n_5916, n6360);
  and g11636 (n6361, n731, n_5916);
  not g11637 (n_5917, n6361);
  and g11638 (n6362, n735, n_5917);
  not g11639 (n_5918, n6362);
  and g11640 (n6363, n739, n_5918);
  not g11641 (n_5919, n6363);
  and g11642 (n6364, n743, n_5919);
  not g11643 (n_5920, n6364);
  and g11644 (n6365, n747, n_5920);
  not g11645 (n_5921, n6365);
  and g11646 (n6366, n751, n_5921);
  not g11647 (n_5922, n6366);
  and g11648 (n6367, n755, n_5922);
  not g11649 (n_5923, n6367);
  and g11650 (n6368, n759, n_5923);
  not g11651 (n_5924, n6368);
  and g11652 (n6369, n763, n_5924);
  not g11653 (n_5925, n6369);
  and g11654 (n6370, n767, n_5925);
  not g11655 (n_5926, n6370);
  and g11656 (n6371, n771, n_5926);
  not g11657 (n_5927, n6371);
  and g11658 (n6372, n775, n_5927);
  not g11659 (n_5928, n6372);
  and g11660 (n6373, n779, n_5928);
  not g11661 (n_5929, n6373);
  and g11662 (n6374, n783, n_5929);
  not g11663 (n_5930, n6374);
  and g11664 (n6375, n787, n_5930);
  not g11665 (n_5931, n6375);
  and g11666 (n6376, n791, n_5931);
  not g11667 (n_5932, n6376);
  and g11668 (n6377, n795, n_5932);
  not g11669 (n_5933, n6377);
  and g11670 (n6378, n799, n_5933);
  not g11671 (n_5934, n6378);
  and g11672 (n6379, n803, n_5934);
  not g11673 (n_5935, n6379);
  and g11674 (n6380, n807, n_5935);
  not g11675 (n_5936, n6380);
  and g11676 (n6381, n811, n_5936);
  not g11677 (n_5937, n6381);
  and g11678 (n6382, n815, n_5937);
  not g11679 (n_5938, n6382);
  and g11680 (n6383, n819, n_5938);
  not g11681 (n_5939, n6383);
  and g11682 (n6384, n823, n_5939);
  not g11683 (n_5940, n6384);
  and g11684 (n6385, n827, n_5940);
  not g11685 (n_5941, n6385);
  and g11686 (n6386, n831, n_5941);
  not g11687 (n_5942, n6386);
  and g11688 (n6387, n835, n_5942);
  not g11689 (n_5943, n6387);
  and g11690 (n6388, n839, n_5943);
  not g11691 (n_5944, n6388);
  and g11692 (n6389, n843, n_5944);
  not g11693 (n_5945, n6389);
  and g11694 (n6390, n847, n_5945);
  not g11695 (n_5946, n6390);
  and g11696 (n6391, n851, n_5946);
  not g11697 (n_5947, n6391);
  and g11698 (n6392, n855, n_5947);
  not g11699 (n_5948, n6392);
  and g11700 (n6393, n859, n_5948);
  not g11701 (n_5949, n6393);
  and g11702 (n6394, n863, n_5949);
  not g11703 (n_5950, n6394);
  and g11704 (n6395, n867, n_5950);
  not g11705 (n_5951, n6395);
  and g11706 (n6396, n871, n_5951);
  not g11707 (n_5952, n6396);
  and g11708 (n6397, n875, n_5952);
  and g11709 (n6398, \req[60] , n_713);
  not g11710 (n_5953, n6397);
  and g11711 (\grant[60] , n_5953, n6398);
  not g11712 (n_5954, n1219);
  and g11713 (n6400, n886, n_5954);
  not g11714 (n_5955, n6400);
  and g11715 (n6401, n891, n_5955);
  not g11716 (n_5956, n6401);
  and g11717 (n6402, n895, n_5956);
  not g11718 (n_5957, n6402);
  and g11719 (n6403, n899, n_5957);
  not g11720 (n_5958, n6403);
  and g11721 (n6404, n903, n_5958);
  not g11722 (n_5959, n6404);
  and g11723 (n6405, n907, n_5959);
  not g11724 (n_5960, n6405);
  and g11725 (n6406, n911, n_5960);
  not g11726 (n_5961, n6406);
  and g11727 (n6407, n915, n_5961);
  not g11728 (n_5962, n6407);
  and g11729 (n6408, n919, n_5962);
  not g11730 (n_5963, n6408);
  and g11731 (n6409, n923, n_5963);
  not g11732 (n_5964, n6409);
  and g11733 (n6410, n927, n_5964);
  not g11734 (n_5965, n6410);
  and g11735 (n6411, n931, n_5965);
  not g11736 (n_5966, n6411);
  and g11737 (n6412, n935, n_5966);
  not g11738 (n_5967, n6412);
  and g11739 (n6413, n939, n_5967);
  not g11740 (n_5968, n6413);
  and g11741 (n6414, n943, n_5968);
  not g11742 (n_5969, n6414);
  and g11743 (n6415, n947, n_5969);
  not g11744 (n_5970, n6415);
  and g11745 (n6416, n951, n_5970);
  not g11746 (n_5971, n6416);
  and g11747 (n6417, n955, n_5971);
  not g11748 (n_5972, n6417);
  and g11749 (n6418, n959, n_5972);
  not g11750 (n_5973, n6418);
  and g11751 (n6419, n963, n_5973);
  not g11752 (n_5974, n6419);
  and g11753 (n6420, n967, n_5974);
  not g11754 (n_5975, n6420);
  and g11755 (n6421, n971, n_5975);
  not g11756 (n_5976, n6421);
  and g11757 (n6422, n975, n_5976);
  not g11758 (n_5977, n6422);
  and g11759 (n6423, n979, n_5977);
  not g11760 (n_5978, n6423);
  and g11761 (n6424, n983, n_5978);
  not g11762 (n_5979, n6424);
  and g11763 (n6425, n987, n_5979);
  not g11764 (n_5980, n6425);
  and g11765 (n6426, n991, n_5980);
  not g11766 (n_5981, n6426);
  and g11767 (n6427, n995, n_5981);
  not g11768 (n_5982, n6427);
  and g11769 (n6428, n999, n_5982);
  not g11770 (n_5983, n6428);
  and g11771 (n6429, n1003, n_5983);
  not g11772 (n_5984, n6429);
  and g11773 (n6430, n1007, n_5984);
  not g11774 (n_5985, n6430);
  and g11775 (n6431, n1011, n_5985);
  not g11776 (n_5986, n6431);
  and g11777 (n6432, n1015, n_5986);
  not g11778 (n_5987, n6432);
  and g11779 (n6433, n1019, n_5987);
  not g11780 (n_5988, n6433);
  and g11781 (n6434, n1023, n_5988);
  not g11782 (n_5989, n6434);
  and g11783 (n6435, n1027, n_5989);
  not g11784 (n_5990, n6435);
  and g11785 (n6436, n1031, n_5990);
  not g11786 (n_5991, n6436);
  and g11787 (n6437, n1035, n_5991);
  not g11788 (n_5992, n6437);
  and g11789 (n6438, n1039, n_5992);
  not g11790 (n_5993, n6438);
  and g11791 (n6439, n1043, n_5993);
  not g11792 (n_5994, n6439);
  and g11793 (n6440, n1047, n_5994);
  not g11794 (n_5995, n6440);
  and g11795 (n6441, n1051, n_5995);
  not g11796 (n_5996, n6441);
  and g11797 (n6442, n1055, n_5996);
  not g11798 (n_5997, n6442);
  and g11799 (n6443, n1059, n_5997);
  not g11800 (n_5998, n6443);
  and g11801 (n6444, n1574, n_5998);
  not g11802 (n_5999, n6444);
  and g11803 (n6445, n1576, n_5999);
  not g11804 (n_6000, n6445);
  and g11805 (n6446, n1837, n_6000);
  not g11806 (n_6001, n6446);
  and g11807 (n6447, n1068, n_6001);
  not g11808 (n_6002, n6447);
  and g11809 (n6448, n1072, n_6002);
  not g11810 (n_6003, n6448);
  and g11811 (n6449, n1076, n_6003);
  not g11812 (n_6004, n6449);
  and g11813 (n6450, n1080, n_6004);
  not g11814 (n_6005, n6450);
  and g11815 (n6451, n1084, n_6005);
  not g11816 (n_6006, n6451);
  and g11817 (n6452, n1088, n_6006);
  not g11818 (n_6007, n6452);
  and g11819 (n6453, n1092, n_6007);
  not g11820 (n_6008, n6453);
  and g11821 (n6454, n1096, n_6008);
  not g11822 (n_6009, n6454);
  and g11823 (n6455, n1100, n_6009);
  not g11824 (n_6010, n6455);
  and g11825 (n6456, n1104, n_6010);
  not g11826 (n_6011, n6456);
  and g11827 (n6457, n1108, n_6011);
  not g11828 (n_6012, n6457);
  and g11829 (n6458, n1112, n_6012);
  not g11830 (n_6013, n6458);
  and g11831 (n6459, n1116, n_6013);
  not g11832 (n_6014, n6459);
  and g11833 (n6460, n1120, n_6014);
  not g11834 (n_6015, n6460);
  and g11835 (n6461, n1124, n_6015);
  not g11836 (n_6016, n6461);
  and g11837 (n6462, n1128, n_6016);
  not g11838 (n_6017, n6462);
  and g11839 (n6463, n1132, n_6017);
  not g11840 (n_6018, n6463);
  and g11841 (n6464, n1136, n_6018);
  not g11842 (n_6019, n6464);
  and g11843 (n6465, n1140, n_6019);
  not g11844 (n_6020, n6465);
  and g11845 (n6466, n1144, n_6020);
  not g11846 (n_6021, n6466);
  and g11847 (n6467, n1148, n_6021);
  not g11848 (n_6022, n6467);
  and g11849 (n6468, n1152, n_6022);
  not g11850 (n_6023, n6468);
  and g11851 (n6469, n1156, n_6023);
  not g11852 (n_6024, n6469);
  and g11853 (n6470, n1160, n_6024);
  not g11854 (n_6025, n6470);
  and g11855 (n6471, n1164, n_6025);
  not g11856 (n_6026, n6471);
  and g11857 (n6472, n1168, n_6026);
  not g11858 (n_6027, n6472);
  and g11859 (n6473, n1172, n_6027);
  not g11860 (n_6028, n6473);
  and g11861 (n6474, n1176, n_6028);
  not g11862 (n_6029, n6474);
  and g11863 (n6475, n1180, n_6029);
  not g11864 (n_6030, n6475);
  and g11865 (n6476, n1184, n_6030);
  not g11866 (n_6031, n6476);
  and g11867 (n6477, n1188, n_6031);
  not g11868 (n_6032, n6477);
  and g11869 (n6478, n1192, n_6032);
  not g11870 (n_6033, n6478);
  and g11871 (n6479, n1196, n_6033);
  not g11872 (n_6034, n6479);
  and g11873 (n6480, n1200, n_6034);
  not g11874 (n_6035, n6480);
  and g11875 (n6481, n1204, n_6035);
  not g11876 (n_6036, n6481);
  and g11877 (n6482, n1208, n_6036);
  not g11878 (n_6037, n6482);
  and g11879 (n6483, n1212, n_6037);
  and g11880 (n6484, \req[61] , n_927);
  not g11881 (n_6038, n6483);
  and g11882 (\grant[61] , n_6038, n6484);
  not g11883 (n_6039, n551);
  and g11884 (n6486, n_6039, n1223);
  not g11885 (n_6040, n6486);
  and g11886 (n6487, n1228, n_6040);
  not g11887 (n_6041, n6487);
  and g11888 (n6488, n1232, n_6041);
  not g11889 (n_6042, n6488);
  and g11890 (n6489, n1236, n_6042);
  not g11891 (n_6043, n6489);
  and g11892 (n6490, n1240, n_6043);
  not g11893 (n_6044, n6490);
  and g11894 (n6491, n1244, n_6044);
  not g11895 (n_6045, n6491);
  and g11896 (n6492, n1248, n_6045);
  not g11897 (n_6046, n6492);
  and g11898 (n6493, n1252, n_6046);
  not g11899 (n_6047, n6493);
  and g11900 (n6494, n1256, n_6047);
  not g11901 (n_6048, n6494);
  and g11902 (n6495, n1260, n_6048);
  not g11903 (n_6049, n6495);
  and g11904 (n6496, n1264, n_6049);
  not g11905 (n_6050, n6496);
  and g11906 (n6497, n1268, n_6050);
  not g11907 (n_6051, n6497);
  and g11908 (n6498, n1272, n_6051);
  not g11909 (n_6052, n6498);
  and g11910 (n6499, n1276, n_6052);
  not g11911 (n_6053, n6499);
  and g11912 (n6500, n1280, n_6053);
  not g11913 (n_6054, n6500);
  and g11914 (n6501, n1284, n_6054);
  not g11915 (n_6055, n6501);
  and g11916 (n6502, n1288, n_6055);
  not g11917 (n_6056, n6502);
  and g11918 (n6503, n1292, n_6056);
  not g11919 (n_6057, n6503);
  and g11920 (n6504, n1296, n_6057);
  not g11921 (n_6058, n6504);
  and g11922 (n6505, n1300, n_6058);
  not g11923 (n_6059, n6505);
  and g11924 (n6506, n1304, n_6059);
  not g11925 (n_6060, n6506);
  and g11926 (n6507, n1308, n_6060);
  not g11927 (n_6061, n6507);
  and g11928 (n6508, n1312, n_6061);
  not g11929 (n_6062, n6508);
  and g11930 (n6509, n1316, n_6062);
  not g11931 (n_6063, n6509);
  and g11932 (n6510, n1320, n_6063);
  not g11933 (n_6064, n6510);
  and g11934 (n6511, n1324, n_6064);
  not g11935 (n_6065, n6511);
  and g11936 (n6512, n1328, n_6065);
  not g11937 (n_6066, n6512);
  and g11938 (n6513, n1332, n_6066);
  not g11939 (n_6067, n6513);
  and g11940 (n6514, n1336, n_6067);
  not g11941 (n_6068, n6514);
  and g11942 (n6515, n1340, n_6068);
  not g11943 (n_6069, n6515);
  and g11944 (n6516, n1344, n_6069);
  not g11945 (n_6070, n6516);
  and g11946 (n6517, n1348, n_6070);
  not g11947 (n_6071, n6517);
  and g11948 (n6518, n1352, n_6071);
  not g11949 (n_6072, n6518);
  and g11950 (n6519, n1356, n_6072);
  not g11951 (n_6073, n6519);
  and g11952 (n6520, n1360, n_6073);
  not g11953 (n_6074, n6520);
  and g11954 (n6521, n1364, n_6074);
  not g11955 (n_6075, n6521);
  and g11956 (n6522, n1368, n_6075);
  not g11957 (n_6076, n6522);
  and g11958 (n6523, n1372, n_6076);
  not g11959 (n_6077, n6523);
  and g11960 (n6524, n1376, n_6077);
  not g11961 (n_6078, n6524);
  and g11962 (n6525, n1380, n_6078);
  not g11963 (n_6079, n6525);
  and g11964 (n6526, n1384, n_6079);
  not g11965 (n_6080, n6526);
  and g11966 (n6527, n1388, n_6080);
  not g11967 (n_6081, n6527);
  and g11968 (n6528, n1392, n_6081);
  not g11969 (n_6082, n6528);
  and g11970 (n6529, n1396, n_6082);
  not g11971 (n_6083, n6529);
  and g11972 (n6530, n1663, n_6083);
  not g11973 (n_6084, n6530);
  and g11974 (n6531, n392, n_6084);
  not g11975 (n_6085, n6531);
  and g11976 (n6532, n396, n_6085);
  not g11977 (n_6086, n6532);
  and g11978 (n6533, n400, n_6086);
  not g11979 (n_6087, n6533);
  and g11980 (n6534, n404, n_6087);
  not g11981 (n_6088, n6534);
  and g11982 (n6535, n408, n_6088);
  not g11983 (n_6089, n6535);
  and g11984 (n6536, n412, n_6089);
  not g11985 (n_6090, n6536);
  and g11986 (n6537, n416, n_6090);
  not g11987 (n_6091, n6537);
  and g11988 (n6538, n420, n_6091);
  not g11989 (n_6092, n6538);
  and g11990 (n6539, n424, n_6092);
  not g11991 (n_6093, n6539);
  and g11992 (n6540, n428, n_6093);
  not g11993 (n_6094, n6540);
  and g11994 (n6541, n432, n_6094);
  not g11995 (n_6095, n6541);
  and g11996 (n6542, n436, n_6095);
  not g11997 (n_6096, n6542);
  and g11998 (n6543, n440, n_6096);
  not g11999 (n_6097, n6543);
  and g12000 (n6544, n444, n_6097);
  not g12001 (n_6098, n6544);
  and g12002 (n6545, n448, n_6098);
  not g12003 (n_6099, n6545);
  and g12004 (n6546, n452, n_6099);
  not g12005 (n_6100, n6546);
  and g12006 (n6547, n456, n_6100);
  not g12007 (n_6101, n6547);
  and g12008 (n6548, n460, n_6101);
  not g12009 (n_6102, n6548);
  and g12010 (n6549, n464, n_6102);
  not g12011 (n_6103, n6549);
  and g12012 (n6550, n468, n_6103);
  not g12013 (n_6104, n6550);
  and g12014 (n6551, n472, n_6104);
  not g12015 (n_6105, n6551);
  and g12016 (n6552, n476, n_6105);
  not g12017 (n_6106, n6552);
  and g12018 (n6553, n480, n_6106);
  not g12019 (n_6107, n6553);
  and g12020 (n6554, n484, n_6107);
  not g12021 (n_6108, n6554);
  and g12022 (n6555, n488, n_6108);
  not g12023 (n_6109, n6555);
  and g12024 (n6556, n492, n_6109);
  not g12025 (n_6110, n6556);
  and g12026 (n6557, n496, n_6110);
  not g12027 (n_6111, n6557);
  and g12028 (n6558, n500, n_6111);
  not g12029 (n_6112, n6558);
  and g12030 (n6559, n504, n_6112);
  not g12031 (n_6113, n6559);
  and g12032 (n6560, n508, n_6113);
  not g12033 (n_6114, n6560);
  and g12034 (n6561, n512, n_6114);
  not g12035 (n_6115, n6561);
  and g12036 (n6562, n516, n_6115);
  not g12037 (n_6116, n6562);
  and g12038 (n6563, n520, n_6116);
  not g12039 (n_6117, n6563);
  and g12040 (n6564, n524, n_6117);
  not g12041 (n_6118, n6564);
  and g12042 (n6565, n528, n_6118);
  not g12043 (n_6119, n6565);
  and g12044 (n6566, n532, n_6119);
  not g12045 (n_6120, n6566);
  and g12046 (n6567, n536, n_6120);
  not g12047 (n_6121, n6567);
  and g12048 (n6568, n540, n_6121);
  not g12049 (n_6122, n6568);
  and g12050 (n6569, n544, n_6122);
  and g12051 (n6570, \req[62] , n_290);
  not g12052 (n_6123, n6569);
  and g12053 (\grant[62] , n_6123, n6570);
  not g12054 (n_6124, n890);
  and g12055 (n6572, n555, n_6124);
  not g12056 (n_6125, n6572);
  and g12057 (n6573, n560, n_6125);
  not g12058 (n_6126, n6573);
  and g12059 (n6574, n564, n_6126);
  not g12060 (n_6127, n6574);
  and g12061 (n6575, n568, n_6127);
  not g12062 (n_6128, n6575);
  and g12063 (n6576, n572, n_6128);
  not g12064 (n_6129, n6576);
  and g12065 (n6577, n576, n_6129);
  not g12066 (n_6130, n6577);
  and g12067 (n6578, n580, n_6130);
  not g12068 (n_6131, n6578);
  and g12069 (n6579, n584, n_6131);
  not g12070 (n_6132, n6579);
  and g12071 (n6580, n588, n_6132);
  not g12072 (n_6133, n6580);
  and g12073 (n6581, n592, n_6133);
  not g12074 (n_6134, n6581);
  and g12075 (n6582, n596, n_6134);
  not g12076 (n_6135, n6582);
  and g12077 (n6583, n600, n_6135);
  not g12078 (n_6136, n6583);
  and g12079 (n6584, n604, n_6136);
  not g12080 (n_6137, n6584);
  and g12081 (n6585, n608, n_6137);
  not g12082 (n_6138, n6585);
  and g12083 (n6586, n612, n_6138);
  not g12084 (n_6139, n6586);
  and g12085 (n6587, n616, n_6139);
  not g12086 (n_6140, n6587);
  and g12087 (n6588, n620, n_6140);
  not g12088 (n_6141, n6588);
  and g12089 (n6589, n624, n_6141);
  not g12090 (n_6142, n6589);
  and g12091 (n6590, n628, n_6142);
  not g12092 (n_6143, n6590);
  and g12093 (n6591, n632, n_6143);
  not g12094 (n_6144, n6591);
  and g12095 (n6592, n636, n_6144);
  not g12096 (n_6145, n6592);
  and g12097 (n6593, n640, n_6145);
  not g12098 (n_6146, n6593);
  and g12099 (n6594, n644, n_6146);
  not g12100 (n_6147, n6594);
  and g12101 (n6595, n648, n_6147);
  not g12102 (n_6148, n6595);
  and g12103 (n6596, n652, n_6148);
  not g12104 (n_6149, n6596);
  and g12105 (n6597, n656, n_6149);
  not g12106 (n_6150, n6597);
  and g12107 (n6598, n660, n_6150);
  not g12108 (n_6151, n6598);
  and g12109 (n6599, n664, n_6151);
  not g12110 (n_6152, n6599);
  and g12111 (n6600, n668, n_6152);
  not g12112 (n_6153, n6600);
  and g12113 (n6601, n672, n_6153);
  not g12114 (n_6154, n6601);
  and g12115 (n6602, n676, n_6154);
  not g12116 (n_6155, n6602);
  and g12117 (n6603, n680, n_6155);
  not g12118 (n_6156, n6603);
  and g12119 (n6604, n684, n_6156);
  not g12120 (n_6157, n6604);
  and g12121 (n6605, n688, n_6157);
  not g12122 (n_6158, n6605);
  and g12123 (n6606, n692, n_6158);
  not g12124 (n_6159, n6606);
  and g12125 (n6607, n696, n_6159);
  not g12126 (n_6160, n6607);
  and g12127 (n6608, n700, n_6160);
  not g12128 (n_6161, n6608);
  and g12129 (n6609, n704, n_6161);
  not g12130 (n_6162, n6609);
  and g12131 (n6610, n708, n_6162);
  not g12132 (n_6163, n6610);
  and g12133 (n6611, n712, n_6163);
  not g12134 (n_6164, n6611);
  and g12135 (n6612, n716, n_6164);
  not g12136 (n_6165, n6612);
  and g12137 (n6613, n720, n_6165);
  not g12138 (n_6166, n6613);
  and g12139 (n6614, n1484, n_6166);
  not g12140 (n_6167, n6614);
  and g12141 (n6615, n1486, n_6167);
  not g12142 (n_6168, n6615);
  and g12143 (n6616, n1750, n_6168);
  not g12144 (n_6169, n6616);
  and g12145 (n6617, n731, n_6169);
  not g12146 (n_6170, n6617);
  and g12147 (n6618, n735, n_6170);
  not g12148 (n_6171, n6618);
  and g12149 (n6619, n739, n_6171);
  not g12150 (n_6172, n6619);
  and g12151 (n6620, n743, n_6172);
  not g12152 (n_6173, n6620);
  and g12153 (n6621, n747, n_6173);
  not g12154 (n_6174, n6621);
  and g12155 (n6622, n751, n_6174);
  not g12156 (n_6175, n6622);
  and g12157 (n6623, n755, n_6175);
  not g12158 (n_6176, n6623);
  and g12159 (n6624, n759, n_6176);
  not g12160 (n_6177, n6624);
  and g12161 (n6625, n763, n_6177);
  not g12162 (n_6178, n6625);
  and g12163 (n6626, n767, n_6178);
  not g12164 (n_6179, n6626);
  and g12165 (n6627, n771, n_6179);
  not g12166 (n_6180, n6627);
  and g12167 (n6628, n775, n_6180);
  not g12168 (n_6181, n6628);
  and g12169 (n6629, n779, n_6181);
  not g12170 (n_6182, n6629);
  and g12171 (n6630, n783, n_6182);
  not g12172 (n_6183, n6630);
  and g12173 (n6631, n787, n_6183);
  not g12174 (n_6184, n6631);
  and g12175 (n6632, n791, n_6184);
  not g12176 (n_6185, n6632);
  and g12177 (n6633, n795, n_6185);
  not g12178 (n_6186, n6633);
  and g12179 (n6634, n799, n_6186);
  not g12180 (n_6187, n6634);
  and g12181 (n6635, n803, n_6187);
  not g12182 (n_6188, n6635);
  and g12183 (n6636, n807, n_6188);
  not g12184 (n_6189, n6636);
  and g12185 (n6637, n811, n_6189);
  not g12186 (n_6190, n6637);
  and g12187 (n6638, n815, n_6190);
  not g12188 (n_6191, n6638);
  and g12189 (n6639, n819, n_6191);
  not g12190 (n_6192, n6639);
  and g12191 (n6640, n823, n_6192);
  not g12192 (n_6193, n6640);
  and g12193 (n6641, n827, n_6193);
  not g12194 (n_6194, n6641);
  and g12195 (n6642, n831, n_6194);
  not g12196 (n_6195, n6642);
  and g12197 (n6643, n835, n_6195);
  not g12198 (n_6196, n6643);
  and g12199 (n6644, n839, n_6196);
  not g12200 (n_6197, n6644);
  and g12201 (n6645, n843, n_6197);
  not g12202 (n_6198, n6645);
  and g12203 (n6646, n847, n_6198);
  not g12204 (n_6199, n6646);
  and g12205 (n6647, n851, n_6199);
  not g12206 (n_6200, n6647);
  and g12207 (n6648, n855, n_6200);
  not g12208 (n_6201, n6648);
  and g12209 (n6649, n859, n_6201);
  not g12210 (n_6202, n6649);
  and g12211 (n6650, n863, n_6202);
  not g12212 (n_6203, n6650);
  and g12213 (n6651, n867, n_6203);
  not g12214 (n_6204, n6651);
  and g12215 (n6652, n871, n_6204);
  not g12216 (n_6205, n6652);
  and g12217 (n6653, n875, n_6205);
  not g12218 (n_6206, n6653);
  and g12219 (n6654, n879, n_6206);
  not g12220 (n_6207, n6654);
  and g12221 (n6655, n883, n_6207);
  and g12222 (n6656, \req[63] , n_719);
  not g12223 (n_6208, n6655);
  and g12224 (\grant[63] , n_6208, n6656);
  not g12225 (n_6209, n1227);
  and g12226 (n6658, n894, n_6209);
  not g12227 (n_6210, n6658);
  and g12228 (n6659, n899, n_6210);
  not g12229 (n_6211, n6659);
  and g12230 (n6660, n903, n_6211);
  not g12231 (n_6212, n6660);
  and g12232 (n6661, n907, n_6212);
  not g12233 (n_6213, n6661);
  and g12234 (n6662, n911, n_6213);
  not g12235 (n_6214, n6662);
  and g12236 (n6663, n915, n_6214);
  not g12237 (n_6215, n6663);
  and g12238 (n6664, n919, n_6215);
  not g12239 (n_6216, n6664);
  and g12240 (n6665, n923, n_6216);
  not g12241 (n_6217, n6665);
  and g12242 (n6666, n927, n_6217);
  not g12243 (n_6218, n6666);
  and g12244 (n6667, n931, n_6218);
  not g12245 (n_6219, n6667);
  and g12246 (n6668, n935, n_6219);
  not g12247 (n_6220, n6668);
  and g12248 (n6669, n939, n_6220);
  not g12249 (n_6221, n6669);
  and g12250 (n6670, n943, n_6221);
  not g12251 (n_6222, n6670);
  and g12252 (n6671, n947, n_6222);
  not g12253 (n_6223, n6671);
  and g12254 (n6672, n951, n_6223);
  not g12255 (n_6224, n6672);
  and g12256 (n6673, n955, n_6224);
  not g12257 (n_6225, n6673);
  and g12258 (n6674, n959, n_6225);
  not g12259 (n_6226, n6674);
  and g12260 (n6675, n963, n_6226);
  not g12261 (n_6227, n6675);
  and g12262 (n6676, n967, n_6227);
  not g12263 (n_6228, n6676);
  and g12264 (n6677, n971, n_6228);
  not g12265 (n_6229, n6677);
  and g12266 (n6678, n975, n_6229);
  not g12267 (n_6230, n6678);
  and g12268 (n6679, n979, n_6230);
  not g12269 (n_6231, n6679);
  and g12270 (n6680, n983, n_6231);
  not g12271 (n_6232, n6680);
  and g12272 (n6681, n987, n_6232);
  not g12273 (n_6233, n6681);
  and g12274 (n6682, n991, n_6233);
  not g12275 (n_6234, n6682);
  and g12276 (n6683, n995, n_6234);
  not g12277 (n_6235, n6683);
  and g12278 (n6684, n999, n_6235);
  not g12279 (n_6236, n6684);
  and g12280 (n6685, n1003, n_6236);
  not g12281 (n_6237, n6685);
  and g12282 (n6686, n1007, n_6237);
  not g12283 (n_6238, n6686);
  and g12284 (n6687, n1011, n_6238);
  not g12285 (n_6239, n6687);
  and g12286 (n6688, n1015, n_6239);
  not g12287 (n_6240, n6688);
  and g12288 (n6689, n1019, n_6240);
  not g12289 (n_6241, n6689);
  and g12290 (n6690, n1023, n_6241);
  not g12291 (n_6242, n6690);
  and g12292 (n6691, n1027, n_6242);
  not g12293 (n_6243, n6691);
  and g12294 (n6692, n1031, n_6243);
  not g12295 (n_6244, n6692);
  and g12296 (n6693, n1035, n_6244);
  not g12297 (n_6245, n6693);
  and g12298 (n6694, n1039, n_6245);
  not g12299 (n_6246, n6694);
  and g12300 (n6695, n1043, n_6246);
  not g12301 (n_6247, n6695);
  and g12302 (n6696, n1047, n_6247);
  not g12303 (n_6248, n6696);
  and g12304 (n6697, n1051, n_6248);
  not g12305 (n_6249, n6697);
  and g12306 (n6698, n1055, n_6249);
  not g12307 (n_6250, n6698);
  and g12308 (n6699, n1059, n_6250);
  not g12309 (n_6251, n6699);
  and g12310 (n6700, n1574, n_6251);
  not g12311 (n_6252, n6700);
  and g12312 (n6701, n1576, n_6252);
  not g12313 (n_6253, n6701);
  and g12314 (n6702, n1837, n_6253);
  not g12315 (n_6254, n6702);
  and g12316 (n6703, n1068, n_6254);
  not g12317 (n_6255, n6703);
  and g12318 (n6704, n1072, n_6255);
  not g12319 (n_6256, n6704);
  and g12320 (n6705, n1076, n_6256);
  not g12321 (n_6257, n6705);
  and g12322 (n6706, n1080, n_6257);
  not g12323 (n_6258, n6706);
  and g12324 (n6707, n1084, n_6258);
  not g12325 (n_6259, n6707);
  and g12326 (n6708, n1088, n_6259);
  not g12327 (n_6260, n6708);
  and g12328 (n6709, n1092, n_6260);
  not g12329 (n_6261, n6709);
  and g12330 (n6710, n1096, n_6261);
  not g12331 (n_6262, n6710);
  and g12332 (n6711, n1100, n_6262);
  not g12333 (n_6263, n6711);
  and g12334 (n6712, n1104, n_6263);
  not g12335 (n_6264, n6712);
  and g12336 (n6713, n1108, n_6264);
  not g12337 (n_6265, n6713);
  and g12338 (n6714, n1112, n_6265);
  not g12339 (n_6266, n6714);
  and g12340 (n6715, n1116, n_6266);
  not g12341 (n_6267, n6715);
  and g12342 (n6716, n1120, n_6267);
  not g12343 (n_6268, n6716);
  and g12344 (n6717, n1124, n_6268);
  not g12345 (n_6269, n6717);
  and g12346 (n6718, n1128, n_6269);
  not g12347 (n_6270, n6718);
  and g12348 (n6719, n1132, n_6270);
  not g12349 (n_6271, n6719);
  and g12350 (n6720, n1136, n_6271);
  not g12351 (n_6272, n6720);
  and g12352 (n6721, n1140, n_6272);
  not g12353 (n_6273, n6721);
  and g12354 (n6722, n1144, n_6273);
  not g12355 (n_6274, n6722);
  and g12356 (n6723, n1148, n_6274);
  not g12357 (n_6275, n6723);
  and g12358 (n6724, n1152, n_6275);
  not g12359 (n_6276, n6724);
  and g12360 (n6725, n1156, n_6276);
  not g12361 (n_6277, n6725);
  and g12362 (n6726, n1160, n_6277);
  not g12363 (n_6278, n6726);
  and g12364 (n6727, n1164, n_6278);
  not g12365 (n_6279, n6727);
  and g12366 (n6728, n1168, n_6279);
  not g12367 (n_6280, n6728);
  and g12368 (n6729, n1172, n_6280);
  not g12369 (n_6281, n6729);
  and g12370 (n6730, n1176, n_6281);
  not g12371 (n_6282, n6730);
  and g12372 (n6731, n1180, n_6282);
  not g12373 (n_6283, n6731);
  and g12374 (n6732, n1184, n_6283);
  not g12375 (n_6284, n6732);
  and g12376 (n6733, n1188, n_6284);
  not g12377 (n_6285, n6733);
  and g12378 (n6734, n1192, n_6285);
  not g12379 (n_6286, n6734);
  and g12380 (n6735, n1196, n_6286);
  not g12381 (n_6287, n6735);
  and g12382 (n6736, n1200, n_6287);
  not g12383 (n_6288, n6736);
  and g12384 (n6737, n1204, n_6288);
  not g12385 (n_6289, n6737);
  and g12386 (n6738, n1208, n_6289);
  not g12387 (n_6290, n6738);
  and g12388 (n6739, n1212, n_6290);
  not g12389 (n_6291, n6739);
  and g12390 (n6740, n1216, n_6291);
  not g12391 (n_6292, n6740);
  and g12392 (n6741, n1220, n_6292);
  and g12393 (n6742, \req[64] , n_931);
  not g12394 (n_6293, n6741);
  and g12395 (\grant[64] , n_6293, n6742);
  not g12396 (n_6294, n559);
  and g12397 (n6744, n_6294, n1231);
  not g12398 (n_6295, n6744);
  and g12399 (n6745, n1236, n_6295);
  not g12400 (n_6296, n6745);
  and g12401 (n6746, n1240, n_6296);
  not g12402 (n_6297, n6746);
  and g12403 (n6747, n1244, n_6297);
  not g12404 (n_6298, n6747);
  and g12405 (n6748, n1248, n_6298);
  not g12406 (n_6299, n6748);
  and g12407 (n6749, n1252, n_6299);
  not g12408 (n_6300, n6749);
  and g12409 (n6750, n1256, n_6300);
  not g12410 (n_6301, n6750);
  and g12411 (n6751, n1260, n_6301);
  not g12412 (n_6302, n6751);
  and g12413 (n6752, n1264, n_6302);
  not g12414 (n_6303, n6752);
  and g12415 (n6753, n1268, n_6303);
  not g12416 (n_6304, n6753);
  and g12417 (n6754, n1272, n_6304);
  not g12418 (n_6305, n6754);
  and g12419 (n6755, n1276, n_6305);
  not g12420 (n_6306, n6755);
  and g12421 (n6756, n1280, n_6306);
  not g12422 (n_6307, n6756);
  and g12423 (n6757, n1284, n_6307);
  not g12424 (n_6308, n6757);
  and g12425 (n6758, n1288, n_6308);
  not g12426 (n_6309, n6758);
  and g12427 (n6759, n1292, n_6309);
  not g12428 (n_6310, n6759);
  and g12429 (n6760, n1296, n_6310);
  not g12430 (n_6311, n6760);
  and g12431 (n6761, n1300, n_6311);
  not g12432 (n_6312, n6761);
  and g12433 (n6762, n1304, n_6312);
  not g12434 (n_6313, n6762);
  and g12435 (n6763, n1308, n_6313);
  not g12436 (n_6314, n6763);
  and g12437 (n6764, n1312, n_6314);
  not g12438 (n_6315, n6764);
  and g12439 (n6765, n1316, n_6315);
  not g12440 (n_6316, n6765);
  and g12441 (n6766, n1320, n_6316);
  not g12442 (n_6317, n6766);
  and g12443 (n6767, n1324, n_6317);
  not g12444 (n_6318, n6767);
  and g12445 (n6768, n1328, n_6318);
  not g12446 (n_6319, n6768);
  and g12447 (n6769, n1332, n_6319);
  not g12448 (n_6320, n6769);
  and g12449 (n6770, n1336, n_6320);
  not g12450 (n_6321, n6770);
  and g12451 (n6771, n1340, n_6321);
  not g12452 (n_6322, n6771);
  and g12453 (n6772, n1344, n_6322);
  not g12454 (n_6323, n6772);
  and g12455 (n6773, n1348, n_6323);
  not g12456 (n_6324, n6773);
  and g12457 (n6774, n1352, n_6324);
  not g12458 (n_6325, n6774);
  and g12459 (n6775, n1356, n_6325);
  not g12460 (n_6326, n6775);
  and g12461 (n6776, n1360, n_6326);
  not g12462 (n_6327, n6776);
  and g12463 (n6777, n1364, n_6327);
  not g12464 (n_6328, n6777);
  and g12465 (n6778, n1368, n_6328);
  not g12466 (n_6329, n6778);
  and g12467 (n6779, n1372, n_6329);
  not g12468 (n_6330, n6779);
  and g12469 (n6780, n1376, n_6330);
  not g12470 (n_6331, n6780);
  and g12471 (n6781, n1380, n_6331);
  not g12472 (n_6332, n6781);
  and g12473 (n6782, n1384, n_6332);
  not g12474 (n_6333, n6782);
  and g12475 (n6783, n1388, n_6333);
  not g12476 (n_6334, n6783);
  and g12477 (n6784, n1392, n_6334);
  not g12478 (n_6335, n6784);
  and g12479 (n6785, n1396, n_6335);
  not g12480 (n_6336, n6785);
  and g12481 (n6786, n1663, n_6336);
  not g12482 (n_6337, n6786);
  and g12483 (n6787, n392, n_6337);
  not g12484 (n_6338, n6787);
  and g12485 (n6788, n396, n_6338);
  not g12486 (n_6339, n6788);
  and g12487 (n6789, n400, n_6339);
  not g12488 (n_6340, n6789);
  and g12489 (n6790, n404, n_6340);
  not g12490 (n_6341, n6790);
  and g12491 (n6791, n408, n_6341);
  not g12492 (n_6342, n6791);
  and g12493 (n6792, n412, n_6342);
  not g12494 (n_6343, n6792);
  and g12495 (n6793, n416, n_6343);
  not g12496 (n_6344, n6793);
  and g12497 (n6794, n420, n_6344);
  not g12498 (n_6345, n6794);
  and g12499 (n6795, n424, n_6345);
  not g12500 (n_6346, n6795);
  and g12501 (n6796, n428, n_6346);
  not g12502 (n_6347, n6796);
  and g12503 (n6797, n432, n_6347);
  not g12504 (n_6348, n6797);
  and g12505 (n6798, n436, n_6348);
  not g12506 (n_6349, n6798);
  and g12507 (n6799, n440, n_6349);
  not g12508 (n_6350, n6799);
  and g12509 (n6800, n444, n_6350);
  not g12510 (n_6351, n6800);
  and g12511 (n6801, n448, n_6351);
  not g12512 (n_6352, n6801);
  and g12513 (n6802, n452, n_6352);
  not g12514 (n_6353, n6802);
  and g12515 (n6803, n456, n_6353);
  not g12516 (n_6354, n6803);
  and g12517 (n6804, n460, n_6354);
  not g12518 (n_6355, n6804);
  and g12519 (n6805, n464, n_6355);
  not g12520 (n_6356, n6805);
  and g12521 (n6806, n468, n_6356);
  not g12522 (n_6357, n6806);
  and g12523 (n6807, n472, n_6357);
  not g12524 (n_6358, n6807);
  and g12525 (n6808, n476, n_6358);
  not g12526 (n_6359, n6808);
  and g12527 (n6809, n480, n_6359);
  not g12528 (n_6360, n6809);
  and g12529 (n6810, n484, n_6360);
  not g12530 (n_6361, n6810);
  and g12531 (n6811, n488, n_6361);
  not g12532 (n_6362, n6811);
  and g12533 (n6812, n492, n_6362);
  not g12534 (n_6363, n6812);
  and g12535 (n6813, n496, n_6363);
  not g12536 (n_6364, n6813);
  and g12537 (n6814, n500, n_6364);
  not g12538 (n_6365, n6814);
  and g12539 (n6815, n504, n_6365);
  not g12540 (n_6366, n6815);
  and g12541 (n6816, n508, n_6366);
  not g12542 (n_6367, n6816);
  and g12543 (n6817, n512, n_6367);
  not g12544 (n_6368, n6817);
  and g12545 (n6818, n516, n_6368);
  not g12546 (n_6369, n6818);
  and g12547 (n6819, n520, n_6369);
  not g12548 (n_6370, n6819);
  and g12549 (n6820, n524, n_6370);
  not g12550 (n_6371, n6820);
  and g12551 (n6821, n528, n_6371);
  not g12552 (n_6372, n6821);
  and g12553 (n6822, n532, n_6372);
  not g12554 (n_6373, n6822);
  and g12555 (n6823, n536, n_6373);
  not g12556 (n_6374, n6823);
  and g12557 (n6824, n540, n_6374);
  not g12558 (n_6375, n6824);
  and g12559 (n6825, n544, n_6375);
  not g12560 (n_6376, n6825);
  and g12561 (n6826, n548, n_6376);
  not g12562 (n_6377, n6826);
  and g12563 (n6827, n552, n_6377);
  and g12564 (n6828, \req[65] , n_304);
  not g12565 (n_6378, n6827);
  and g12566 (\grant[65] , n_6378, n6828);
  not g12567 (n_6379, n898);
  and g12568 (n6830, n563, n_6379);
  not g12569 (n_6380, n6830);
  and g12570 (n6831, n568, n_6380);
  not g12571 (n_6381, n6831);
  and g12572 (n6832, n572, n_6381);
  not g12573 (n_6382, n6832);
  and g12574 (n6833, n576, n_6382);
  not g12575 (n_6383, n6833);
  and g12576 (n6834, n580, n_6383);
  not g12577 (n_6384, n6834);
  and g12578 (n6835, n584, n_6384);
  not g12579 (n_6385, n6835);
  and g12580 (n6836, n588, n_6385);
  not g12581 (n_6386, n6836);
  and g12582 (n6837, n592, n_6386);
  not g12583 (n_6387, n6837);
  and g12584 (n6838, n596, n_6387);
  not g12585 (n_6388, n6838);
  and g12586 (n6839, n600, n_6388);
  not g12587 (n_6389, n6839);
  and g12588 (n6840, n604, n_6389);
  not g12589 (n_6390, n6840);
  and g12590 (n6841, n608, n_6390);
  not g12591 (n_6391, n6841);
  and g12592 (n6842, n612, n_6391);
  not g12593 (n_6392, n6842);
  and g12594 (n6843, n616, n_6392);
  not g12595 (n_6393, n6843);
  and g12596 (n6844, n620, n_6393);
  not g12597 (n_6394, n6844);
  and g12598 (n6845, n624, n_6394);
  not g12599 (n_6395, n6845);
  and g12600 (n6846, n628, n_6395);
  not g12601 (n_6396, n6846);
  and g12602 (n6847, n632, n_6396);
  not g12603 (n_6397, n6847);
  and g12604 (n6848, n636, n_6397);
  not g12605 (n_6398, n6848);
  and g12606 (n6849, n640, n_6398);
  not g12607 (n_6399, n6849);
  and g12608 (n6850, n644, n_6399);
  not g12609 (n_6400, n6850);
  and g12610 (n6851, n648, n_6400);
  not g12611 (n_6401, n6851);
  and g12612 (n6852, n652, n_6401);
  not g12613 (n_6402, n6852);
  and g12614 (n6853, n656, n_6402);
  not g12615 (n_6403, n6853);
  and g12616 (n6854, n660, n_6403);
  not g12617 (n_6404, n6854);
  and g12618 (n6855, n664, n_6404);
  not g12619 (n_6405, n6855);
  and g12620 (n6856, n668, n_6405);
  not g12621 (n_6406, n6856);
  and g12622 (n6857, n672, n_6406);
  not g12623 (n_6407, n6857);
  and g12624 (n6858, n676, n_6407);
  not g12625 (n_6408, n6858);
  and g12626 (n6859, n680, n_6408);
  not g12627 (n_6409, n6859);
  and g12628 (n6860, n684, n_6409);
  not g12629 (n_6410, n6860);
  and g12630 (n6861, n688, n_6410);
  not g12631 (n_6411, n6861);
  and g12632 (n6862, n692, n_6411);
  not g12633 (n_6412, n6862);
  and g12634 (n6863, n696, n_6412);
  not g12635 (n_6413, n6863);
  and g12636 (n6864, n700, n_6413);
  not g12637 (n_6414, n6864);
  and g12638 (n6865, n704, n_6414);
  not g12639 (n_6415, n6865);
  and g12640 (n6866, n708, n_6415);
  not g12641 (n_6416, n6866);
  and g12642 (n6867, n712, n_6416);
  not g12643 (n_6417, n6867);
  and g12644 (n6868, n716, n_6417);
  not g12645 (n_6418, n6868);
  and g12646 (n6869, n720, n_6418);
  not g12647 (n_6419, n6869);
  and g12648 (n6870, n1484, n_6419);
  not g12649 (n_6420, n6870);
  and g12650 (n6871, n1486, n_6420);
  not g12651 (n_6421, n6871);
  and g12652 (n6872, n1750, n_6421);
  not g12653 (n_6422, n6872);
  and g12654 (n6873, n731, n_6422);
  not g12655 (n_6423, n6873);
  and g12656 (n6874, n735, n_6423);
  not g12657 (n_6424, n6874);
  and g12658 (n6875, n739, n_6424);
  not g12659 (n_6425, n6875);
  and g12660 (n6876, n743, n_6425);
  not g12661 (n_6426, n6876);
  and g12662 (n6877, n747, n_6426);
  not g12663 (n_6427, n6877);
  and g12664 (n6878, n751, n_6427);
  not g12665 (n_6428, n6878);
  and g12666 (n6879, n755, n_6428);
  not g12667 (n_6429, n6879);
  and g12668 (n6880, n759, n_6429);
  not g12669 (n_6430, n6880);
  and g12670 (n6881, n763, n_6430);
  not g12671 (n_6431, n6881);
  and g12672 (n6882, n767, n_6431);
  not g12673 (n_6432, n6882);
  and g12674 (n6883, n771, n_6432);
  not g12675 (n_6433, n6883);
  and g12676 (n6884, n775, n_6433);
  not g12677 (n_6434, n6884);
  and g12678 (n6885, n779, n_6434);
  not g12679 (n_6435, n6885);
  and g12680 (n6886, n783, n_6435);
  not g12681 (n_6436, n6886);
  and g12682 (n6887, n787, n_6436);
  not g12683 (n_6437, n6887);
  and g12684 (n6888, n791, n_6437);
  not g12685 (n_6438, n6888);
  and g12686 (n6889, n795, n_6438);
  not g12687 (n_6439, n6889);
  and g12688 (n6890, n799, n_6439);
  not g12689 (n_6440, n6890);
  and g12690 (n6891, n803, n_6440);
  not g12691 (n_6441, n6891);
  and g12692 (n6892, n807, n_6441);
  not g12693 (n_6442, n6892);
  and g12694 (n6893, n811, n_6442);
  not g12695 (n_6443, n6893);
  and g12696 (n6894, n815, n_6443);
  not g12697 (n_6444, n6894);
  and g12698 (n6895, n819, n_6444);
  not g12699 (n_6445, n6895);
  and g12700 (n6896, n823, n_6445);
  not g12701 (n_6446, n6896);
  and g12702 (n6897, n827, n_6446);
  not g12703 (n_6447, n6897);
  and g12704 (n6898, n831, n_6447);
  not g12705 (n_6448, n6898);
  and g12706 (n6899, n835, n_6448);
  not g12707 (n_6449, n6899);
  and g12708 (n6900, n839, n_6449);
  not g12709 (n_6450, n6900);
  and g12710 (n6901, n843, n_6450);
  not g12711 (n_6451, n6901);
  and g12712 (n6902, n847, n_6451);
  not g12713 (n_6452, n6902);
  and g12714 (n6903, n851, n_6452);
  not g12715 (n_6453, n6903);
  and g12716 (n6904, n855, n_6453);
  not g12717 (n_6454, n6904);
  and g12718 (n6905, n859, n_6454);
  not g12719 (n_6455, n6905);
  and g12720 (n6906, n863, n_6455);
  not g12721 (n_6456, n6906);
  and g12722 (n6907, n867, n_6456);
  not g12723 (n_6457, n6907);
  and g12724 (n6908, n871, n_6457);
  not g12725 (n_6458, n6908);
  and g12726 (n6909, n875, n_6458);
  not g12727 (n_6459, n6909);
  and g12728 (n6910, n879, n_6459);
  not g12729 (n_6460, n6910);
  and g12730 (n6911, n883, n_6460);
  not g12731 (n_6461, n6911);
  and g12732 (n6912, n887, n_6461);
  not g12733 (n_6462, n6912);
  and g12734 (n6913, n891, n_6462);
  and g12735 (n6914, \req[66] , n_725);
  not g12736 (n_6463, n6913);
  and g12737 (\grant[66] , n_6463, n6914);
  not g12738 (n_6464, n1235);
  and g12739 (n6916, n902, n_6464);
  not g12740 (n_6465, n6916);
  and g12741 (n6917, n907, n_6465);
  not g12742 (n_6466, n6917);
  and g12743 (n6918, n911, n_6466);
  not g12744 (n_6467, n6918);
  and g12745 (n6919, n915, n_6467);
  not g12746 (n_6468, n6919);
  and g12747 (n6920, n919, n_6468);
  not g12748 (n_6469, n6920);
  and g12749 (n6921, n923, n_6469);
  not g12750 (n_6470, n6921);
  and g12751 (n6922, n927, n_6470);
  not g12752 (n_6471, n6922);
  and g12753 (n6923, n931, n_6471);
  not g12754 (n_6472, n6923);
  and g12755 (n6924, n935, n_6472);
  not g12756 (n_6473, n6924);
  and g12757 (n6925, n939, n_6473);
  not g12758 (n_6474, n6925);
  and g12759 (n6926, n943, n_6474);
  not g12760 (n_6475, n6926);
  and g12761 (n6927, n947, n_6475);
  not g12762 (n_6476, n6927);
  and g12763 (n6928, n951, n_6476);
  not g12764 (n_6477, n6928);
  and g12765 (n6929, n955, n_6477);
  not g12766 (n_6478, n6929);
  and g12767 (n6930, n959, n_6478);
  not g12768 (n_6479, n6930);
  and g12769 (n6931, n963, n_6479);
  not g12770 (n_6480, n6931);
  and g12771 (n6932, n967, n_6480);
  not g12772 (n_6481, n6932);
  and g12773 (n6933, n971, n_6481);
  not g12774 (n_6482, n6933);
  and g12775 (n6934, n975, n_6482);
  not g12776 (n_6483, n6934);
  and g12777 (n6935, n979, n_6483);
  not g12778 (n_6484, n6935);
  and g12779 (n6936, n983, n_6484);
  not g12780 (n_6485, n6936);
  and g12781 (n6937, n987, n_6485);
  not g12782 (n_6486, n6937);
  and g12783 (n6938, n991, n_6486);
  not g12784 (n_6487, n6938);
  and g12785 (n6939, n995, n_6487);
  not g12786 (n_6488, n6939);
  and g12787 (n6940, n999, n_6488);
  not g12788 (n_6489, n6940);
  and g12789 (n6941, n1003, n_6489);
  not g12790 (n_6490, n6941);
  and g12791 (n6942, n1007, n_6490);
  not g12792 (n_6491, n6942);
  and g12793 (n6943, n1011, n_6491);
  not g12794 (n_6492, n6943);
  and g12795 (n6944, n1015, n_6492);
  not g12796 (n_6493, n6944);
  and g12797 (n6945, n1019, n_6493);
  not g12798 (n_6494, n6945);
  and g12799 (n6946, n1023, n_6494);
  not g12800 (n_6495, n6946);
  and g12801 (n6947, n1027, n_6495);
  not g12802 (n_6496, n6947);
  and g12803 (n6948, n1031, n_6496);
  not g12804 (n_6497, n6948);
  and g12805 (n6949, n1035, n_6497);
  not g12806 (n_6498, n6949);
  and g12807 (n6950, n1039, n_6498);
  not g12808 (n_6499, n6950);
  and g12809 (n6951, n1043, n_6499);
  not g12810 (n_6500, n6951);
  and g12811 (n6952, n1047, n_6500);
  not g12812 (n_6501, n6952);
  and g12813 (n6953, n1051, n_6501);
  not g12814 (n_6502, n6953);
  and g12815 (n6954, n1055, n_6502);
  not g12816 (n_6503, n6954);
  and g12817 (n6955, n1059, n_6503);
  not g12818 (n_6504, n6955);
  and g12819 (n6956, n1574, n_6504);
  not g12820 (n_6505, n6956);
  and g12821 (n6957, n1576, n_6505);
  not g12822 (n_6506, n6957);
  and g12823 (n6958, n1837, n_6506);
  not g12824 (n_6507, n6958);
  and g12825 (n6959, n1068, n_6507);
  not g12826 (n_6508, n6959);
  and g12827 (n6960, n1072, n_6508);
  not g12828 (n_6509, n6960);
  and g12829 (n6961, n1076, n_6509);
  not g12830 (n_6510, n6961);
  and g12831 (n6962, n1080, n_6510);
  not g12832 (n_6511, n6962);
  and g12833 (n6963, n1084, n_6511);
  not g12834 (n_6512, n6963);
  and g12835 (n6964, n1088, n_6512);
  not g12836 (n_6513, n6964);
  and g12837 (n6965, n1092, n_6513);
  not g12838 (n_6514, n6965);
  and g12839 (n6966, n1096, n_6514);
  not g12840 (n_6515, n6966);
  and g12841 (n6967, n1100, n_6515);
  not g12842 (n_6516, n6967);
  and g12843 (n6968, n1104, n_6516);
  not g12844 (n_6517, n6968);
  and g12845 (n6969, n1108, n_6517);
  not g12846 (n_6518, n6969);
  and g12847 (n6970, n1112, n_6518);
  not g12848 (n_6519, n6970);
  and g12849 (n6971, n1116, n_6519);
  not g12850 (n_6520, n6971);
  and g12851 (n6972, n1120, n_6520);
  not g12852 (n_6521, n6972);
  and g12853 (n6973, n1124, n_6521);
  not g12854 (n_6522, n6973);
  and g12855 (n6974, n1128, n_6522);
  not g12856 (n_6523, n6974);
  and g12857 (n6975, n1132, n_6523);
  not g12858 (n_6524, n6975);
  and g12859 (n6976, n1136, n_6524);
  not g12860 (n_6525, n6976);
  and g12861 (n6977, n1140, n_6525);
  not g12862 (n_6526, n6977);
  and g12863 (n6978, n1144, n_6526);
  not g12864 (n_6527, n6978);
  and g12865 (n6979, n1148, n_6527);
  not g12866 (n_6528, n6979);
  and g12867 (n6980, n1152, n_6528);
  not g12868 (n_6529, n6980);
  and g12869 (n6981, n1156, n_6529);
  not g12870 (n_6530, n6981);
  and g12871 (n6982, n1160, n_6530);
  not g12872 (n_6531, n6982);
  and g12873 (n6983, n1164, n_6531);
  not g12874 (n_6532, n6983);
  and g12875 (n6984, n1168, n_6532);
  not g12876 (n_6533, n6984);
  and g12877 (n6985, n1172, n_6533);
  not g12878 (n_6534, n6985);
  and g12879 (n6986, n1176, n_6534);
  not g12880 (n_6535, n6986);
  and g12881 (n6987, n1180, n_6535);
  not g12882 (n_6536, n6987);
  and g12883 (n6988, n1184, n_6536);
  not g12884 (n_6537, n6988);
  and g12885 (n6989, n1188, n_6537);
  not g12886 (n_6538, n6989);
  and g12887 (n6990, n1192, n_6538);
  not g12888 (n_6539, n6990);
  and g12889 (n6991, n1196, n_6539);
  not g12890 (n_6540, n6991);
  and g12891 (n6992, n1200, n_6540);
  not g12892 (n_6541, n6992);
  and g12893 (n6993, n1204, n_6541);
  not g12894 (n_6542, n6993);
  and g12895 (n6994, n1208, n_6542);
  not g12896 (n_6543, n6994);
  and g12897 (n6995, n1212, n_6543);
  not g12898 (n_6544, n6995);
  and g12899 (n6996, n1216, n_6544);
  not g12900 (n_6545, n6996);
  and g12901 (n6997, n1220, n_6545);
  not g12902 (n_6546, n6997);
  and g12903 (n6998, n1224, n_6546);
  not g12904 (n_6547, n6998);
  and g12905 (n6999, n1228, n_6547);
  and g12906 (n7000, \req[67] , n_935);
  not g12907 (n_6548, n6999);
  and g12908 (\grant[67] , n_6548, n7000);
  not g12909 (n_6549, n567);
  and g12910 (n7002, n_6549, n1239);
  not g12911 (n_6550, n7002);
  and g12912 (n7003, n1244, n_6550);
  not g12913 (n_6551, n7003);
  and g12914 (n7004, n1248, n_6551);
  not g12915 (n_6552, n7004);
  and g12916 (n7005, n1252, n_6552);
  not g12917 (n_6553, n7005);
  and g12918 (n7006, n1256, n_6553);
  not g12919 (n_6554, n7006);
  and g12920 (n7007, n1260, n_6554);
  not g12921 (n_6555, n7007);
  and g12922 (n7008, n1264, n_6555);
  not g12923 (n_6556, n7008);
  and g12924 (n7009, n1268, n_6556);
  not g12925 (n_6557, n7009);
  and g12926 (n7010, n1272, n_6557);
  not g12927 (n_6558, n7010);
  and g12928 (n7011, n1276, n_6558);
  not g12929 (n_6559, n7011);
  and g12930 (n7012, n1280, n_6559);
  not g12931 (n_6560, n7012);
  and g12932 (n7013, n1284, n_6560);
  not g12933 (n_6561, n7013);
  and g12934 (n7014, n1288, n_6561);
  not g12935 (n_6562, n7014);
  and g12936 (n7015, n1292, n_6562);
  not g12937 (n_6563, n7015);
  and g12938 (n7016, n1296, n_6563);
  not g12939 (n_6564, n7016);
  and g12940 (n7017, n1300, n_6564);
  not g12941 (n_6565, n7017);
  and g12942 (n7018, n1304, n_6565);
  not g12943 (n_6566, n7018);
  and g12944 (n7019, n1308, n_6566);
  not g12945 (n_6567, n7019);
  and g12946 (n7020, n1312, n_6567);
  not g12947 (n_6568, n7020);
  and g12948 (n7021, n1316, n_6568);
  not g12949 (n_6569, n7021);
  and g12950 (n7022, n1320, n_6569);
  not g12951 (n_6570, n7022);
  and g12952 (n7023, n1324, n_6570);
  not g12953 (n_6571, n7023);
  and g12954 (n7024, n1328, n_6571);
  not g12955 (n_6572, n7024);
  and g12956 (n7025, n1332, n_6572);
  not g12957 (n_6573, n7025);
  and g12958 (n7026, n1336, n_6573);
  not g12959 (n_6574, n7026);
  and g12960 (n7027, n1340, n_6574);
  not g12961 (n_6575, n7027);
  and g12962 (n7028, n1344, n_6575);
  not g12963 (n_6576, n7028);
  and g12964 (n7029, n1348, n_6576);
  not g12965 (n_6577, n7029);
  and g12966 (n7030, n1352, n_6577);
  not g12967 (n_6578, n7030);
  and g12968 (n7031, n1356, n_6578);
  not g12969 (n_6579, n7031);
  and g12970 (n7032, n1360, n_6579);
  not g12971 (n_6580, n7032);
  and g12972 (n7033, n1364, n_6580);
  not g12973 (n_6581, n7033);
  and g12974 (n7034, n1368, n_6581);
  not g12975 (n_6582, n7034);
  and g12976 (n7035, n1372, n_6582);
  not g12977 (n_6583, n7035);
  and g12978 (n7036, n1376, n_6583);
  not g12979 (n_6584, n7036);
  and g12980 (n7037, n1380, n_6584);
  not g12981 (n_6585, n7037);
  and g12982 (n7038, n1384, n_6585);
  not g12983 (n_6586, n7038);
  and g12984 (n7039, n1388, n_6586);
  not g12985 (n_6587, n7039);
  and g12986 (n7040, n1392, n_6587);
  not g12987 (n_6588, n7040);
  and g12988 (n7041, n1396, n_6588);
  not g12989 (n_6589, n7041);
  and g12990 (n7042, n1663, n_6589);
  not g12991 (n_6590, n7042);
  and g12992 (n7043, n392, n_6590);
  not g12993 (n_6591, n7043);
  and g12994 (n7044, n396, n_6591);
  not g12995 (n_6592, n7044);
  and g12996 (n7045, n400, n_6592);
  not g12997 (n_6593, n7045);
  and g12998 (n7046, n404, n_6593);
  not g12999 (n_6594, n7046);
  and g13000 (n7047, n408, n_6594);
  not g13001 (n_6595, n7047);
  and g13002 (n7048, n412, n_6595);
  not g13003 (n_6596, n7048);
  and g13004 (n7049, n416, n_6596);
  not g13005 (n_6597, n7049);
  and g13006 (n7050, n420, n_6597);
  not g13007 (n_6598, n7050);
  and g13008 (n7051, n424, n_6598);
  not g13009 (n_6599, n7051);
  and g13010 (n7052, n428, n_6599);
  not g13011 (n_6600, n7052);
  and g13012 (n7053, n432, n_6600);
  not g13013 (n_6601, n7053);
  and g13014 (n7054, n436, n_6601);
  not g13015 (n_6602, n7054);
  and g13016 (n7055, n440, n_6602);
  not g13017 (n_6603, n7055);
  and g13018 (n7056, n444, n_6603);
  not g13019 (n_6604, n7056);
  and g13020 (n7057, n448, n_6604);
  not g13021 (n_6605, n7057);
  and g13022 (n7058, n452, n_6605);
  not g13023 (n_6606, n7058);
  and g13024 (n7059, n456, n_6606);
  not g13025 (n_6607, n7059);
  and g13026 (n7060, n460, n_6607);
  not g13027 (n_6608, n7060);
  and g13028 (n7061, n464, n_6608);
  not g13029 (n_6609, n7061);
  and g13030 (n7062, n468, n_6609);
  not g13031 (n_6610, n7062);
  and g13032 (n7063, n472, n_6610);
  not g13033 (n_6611, n7063);
  and g13034 (n7064, n476, n_6611);
  not g13035 (n_6612, n7064);
  and g13036 (n7065, n480, n_6612);
  not g13037 (n_6613, n7065);
  and g13038 (n7066, n484, n_6613);
  not g13039 (n_6614, n7066);
  and g13040 (n7067, n488, n_6614);
  not g13041 (n_6615, n7067);
  and g13042 (n7068, n492, n_6615);
  not g13043 (n_6616, n7068);
  and g13044 (n7069, n496, n_6616);
  not g13045 (n_6617, n7069);
  and g13046 (n7070, n500, n_6617);
  not g13047 (n_6618, n7070);
  and g13048 (n7071, n504, n_6618);
  not g13049 (n_6619, n7071);
  and g13050 (n7072, n508, n_6619);
  not g13051 (n_6620, n7072);
  and g13052 (n7073, n512, n_6620);
  not g13053 (n_6621, n7073);
  and g13054 (n7074, n516, n_6621);
  not g13055 (n_6622, n7074);
  and g13056 (n7075, n520, n_6622);
  not g13057 (n_6623, n7075);
  and g13058 (n7076, n524, n_6623);
  not g13059 (n_6624, n7076);
  and g13060 (n7077, n528, n_6624);
  not g13061 (n_6625, n7077);
  and g13062 (n7078, n532, n_6625);
  not g13063 (n_6626, n7078);
  and g13064 (n7079, n536, n_6626);
  not g13065 (n_6627, n7079);
  and g13066 (n7080, n540, n_6627);
  not g13067 (n_6628, n7080);
  and g13068 (n7081, n544, n_6628);
  not g13069 (n_6629, n7081);
  and g13070 (n7082, n548, n_6629);
  not g13071 (n_6630, n7082);
  and g13072 (n7083, n552, n_6630);
  not g13073 (n_6631, n7083);
  and g13074 (n7084, n556, n_6631);
  not g13075 (n_6632, n7084);
  and g13076 (n7085, n560, n_6632);
  and g13077 (n7086, \req[68] , n_318);
  not g13078 (n_6633, n7085);
  and g13079 (\grant[68] , n_6633, n7086);
  not g13080 (n_6634, n906);
  and g13081 (n7088, n571, n_6634);
  not g13082 (n_6635, n7088);
  and g13083 (n7089, n576, n_6635);
  not g13084 (n_6636, n7089);
  and g13085 (n7090, n580, n_6636);
  not g13086 (n_6637, n7090);
  and g13087 (n7091, n584, n_6637);
  not g13088 (n_6638, n7091);
  and g13089 (n7092, n588, n_6638);
  not g13090 (n_6639, n7092);
  and g13091 (n7093, n592, n_6639);
  not g13092 (n_6640, n7093);
  and g13093 (n7094, n596, n_6640);
  not g13094 (n_6641, n7094);
  and g13095 (n7095, n600, n_6641);
  not g13096 (n_6642, n7095);
  and g13097 (n7096, n604, n_6642);
  not g13098 (n_6643, n7096);
  and g13099 (n7097, n608, n_6643);
  not g13100 (n_6644, n7097);
  and g13101 (n7098, n612, n_6644);
  not g13102 (n_6645, n7098);
  and g13103 (n7099, n616, n_6645);
  not g13104 (n_6646, n7099);
  and g13105 (n7100, n620, n_6646);
  not g13106 (n_6647, n7100);
  and g13107 (n7101, n624, n_6647);
  not g13108 (n_6648, n7101);
  and g13109 (n7102, n628, n_6648);
  not g13110 (n_6649, n7102);
  and g13111 (n7103, n632, n_6649);
  not g13112 (n_6650, n7103);
  and g13113 (n7104, n636, n_6650);
  not g13114 (n_6651, n7104);
  and g13115 (n7105, n640, n_6651);
  not g13116 (n_6652, n7105);
  and g13117 (n7106, n644, n_6652);
  not g13118 (n_6653, n7106);
  and g13119 (n7107, n648, n_6653);
  not g13120 (n_6654, n7107);
  and g13121 (n7108, n652, n_6654);
  not g13122 (n_6655, n7108);
  and g13123 (n7109, n656, n_6655);
  not g13124 (n_6656, n7109);
  and g13125 (n7110, n660, n_6656);
  not g13126 (n_6657, n7110);
  and g13127 (n7111, n664, n_6657);
  not g13128 (n_6658, n7111);
  and g13129 (n7112, n668, n_6658);
  not g13130 (n_6659, n7112);
  and g13131 (n7113, n672, n_6659);
  not g13132 (n_6660, n7113);
  and g13133 (n7114, n676, n_6660);
  not g13134 (n_6661, n7114);
  and g13135 (n7115, n680, n_6661);
  not g13136 (n_6662, n7115);
  and g13137 (n7116, n684, n_6662);
  not g13138 (n_6663, n7116);
  and g13139 (n7117, n688, n_6663);
  not g13140 (n_6664, n7117);
  and g13141 (n7118, n692, n_6664);
  not g13142 (n_6665, n7118);
  and g13143 (n7119, n696, n_6665);
  not g13144 (n_6666, n7119);
  and g13145 (n7120, n700, n_6666);
  not g13146 (n_6667, n7120);
  and g13147 (n7121, n704, n_6667);
  not g13148 (n_6668, n7121);
  and g13149 (n7122, n708, n_6668);
  not g13150 (n_6669, n7122);
  and g13151 (n7123, n712, n_6669);
  not g13152 (n_6670, n7123);
  and g13153 (n7124, n716, n_6670);
  not g13154 (n_6671, n7124);
  and g13155 (n7125, n720, n_6671);
  not g13156 (n_6672, n7125);
  and g13157 (n7126, n1484, n_6672);
  not g13158 (n_6673, n7126);
  and g13159 (n7127, n1486, n_6673);
  not g13160 (n_6674, n7127);
  and g13161 (n7128, n1750, n_6674);
  not g13162 (n_6675, n7128);
  and g13163 (n7129, n731, n_6675);
  not g13164 (n_6676, n7129);
  and g13165 (n7130, n735, n_6676);
  not g13166 (n_6677, n7130);
  and g13167 (n7131, n739, n_6677);
  not g13168 (n_6678, n7131);
  and g13169 (n7132, n743, n_6678);
  not g13170 (n_6679, n7132);
  and g13171 (n7133, n747, n_6679);
  not g13172 (n_6680, n7133);
  and g13173 (n7134, n751, n_6680);
  not g13174 (n_6681, n7134);
  and g13175 (n7135, n755, n_6681);
  not g13176 (n_6682, n7135);
  and g13177 (n7136, n759, n_6682);
  not g13178 (n_6683, n7136);
  and g13179 (n7137, n763, n_6683);
  not g13180 (n_6684, n7137);
  and g13181 (n7138, n767, n_6684);
  not g13182 (n_6685, n7138);
  and g13183 (n7139, n771, n_6685);
  not g13184 (n_6686, n7139);
  and g13185 (n7140, n775, n_6686);
  not g13186 (n_6687, n7140);
  and g13187 (n7141, n779, n_6687);
  not g13188 (n_6688, n7141);
  and g13189 (n7142, n783, n_6688);
  not g13190 (n_6689, n7142);
  and g13191 (n7143, n787, n_6689);
  not g13192 (n_6690, n7143);
  and g13193 (n7144, n791, n_6690);
  not g13194 (n_6691, n7144);
  and g13195 (n7145, n795, n_6691);
  not g13196 (n_6692, n7145);
  and g13197 (n7146, n799, n_6692);
  not g13198 (n_6693, n7146);
  and g13199 (n7147, n803, n_6693);
  not g13200 (n_6694, n7147);
  and g13201 (n7148, n807, n_6694);
  not g13202 (n_6695, n7148);
  and g13203 (n7149, n811, n_6695);
  not g13204 (n_6696, n7149);
  and g13205 (n7150, n815, n_6696);
  not g13206 (n_6697, n7150);
  and g13207 (n7151, n819, n_6697);
  not g13208 (n_6698, n7151);
  and g13209 (n7152, n823, n_6698);
  not g13210 (n_6699, n7152);
  and g13211 (n7153, n827, n_6699);
  not g13212 (n_6700, n7153);
  and g13213 (n7154, n831, n_6700);
  not g13214 (n_6701, n7154);
  and g13215 (n7155, n835, n_6701);
  not g13216 (n_6702, n7155);
  and g13217 (n7156, n839, n_6702);
  not g13218 (n_6703, n7156);
  and g13219 (n7157, n843, n_6703);
  not g13220 (n_6704, n7157);
  and g13221 (n7158, n847, n_6704);
  not g13222 (n_6705, n7158);
  and g13223 (n7159, n851, n_6705);
  not g13224 (n_6706, n7159);
  and g13225 (n7160, n855, n_6706);
  not g13226 (n_6707, n7160);
  and g13227 (n7161, n859, n_6707);
  not g13228 (n_6708, n7161);
  and g13229 (n7162, n863, n_6708);
  not g13230 (n_6709, n7162);
  and g13231 (n7163, n867, n_6709);
  not g13232 (n_6710, n7163);
  and g13233 (n7164, n871, n_6710);
  not g13234 (n_6711, n7164);
  and g13235 (n7165, n875, n_6711);
  not g13236 (n_6712, n7165);
  and g13237 (n7166, n879, n_6712);
  not g13238 (n_6713, n7166);
  and g13239 (n7167, n883, n_6713);
  not g13240 (n_6714, n7167);
  and g13241 (n7168, n887, n_6714);
  not g13242 (n_6715, n7168);
  and g13243 (n7169, n891, n_6715);
  not g13244 (n_6716, n7169);
  and g13245 (n7170, n895, n_6716);
  not g13246 (n_6717, n7170);
  and g13247 (n7171, n899, n_6717);
  and g13248 (n7172, \req[69] , n_731);
  not g13249 (n_6718, n7171);
  and g13250 (\grant[69] , n_6718, n7172);
  not g13251 (n_6719, n1243);
  and g13252 (n7174, n910, n_6719);
  not g13253 (n_6720, n7174);
  and g13254 (n7175, n915, n_6720);
  not g13255 (n_6721, n7175);
  and g13256 (n7176, n919, n_6721);
  not g13257 (n_6722, n7176);
  and g13258 (n7177, n923, n_6722);
  not g13259 (n_6723, n7177);
  and g13260 (n7178, n927, n_6723);
  not g13261 (n_6724, n7178);
  and g13262 (n7179, n931, n_6724);
  not g13263 (n_6725, n7179);
  and g13264 (n7180, n935, n_6725);
  not g13265 (n_6726, n7180);
  and g13266 (n7181, n939, n_6726);
  not g13267 (n_6727, n7181);
  and g13268 (n7182, n943, n_6727);
  not g13269 (n_6728, n7182);
  and g13270 (n7183, n947, n_6728);
  not g13271 (n_6729, n7183);
  and g13272 (n7184, n951, n_6729);
  not g13273 (n_6730, n7184);
  and g13274 (n7185, n955, n_6730);
  not g13275 (n_6731, n7185);
  and g13276 (n7186, n959, n_6731);
  not g13277 (n_6732, n7186);
  and g13278 (n7187, n963, n_6732);
  not g13279 (n_6733, n7187);
  and g13280 (n7188, n967, n_6733);
  not g13281 (n_6734, n7188);
  and g13282 (n7189, n971, n_6734);
  not g13283 (n_6735, n7189);
  and g13284 (n7190, n975, n_6735);
  not g13285 (n_6736, n7190);
  and g13286 (n7191, n979, n_6736);
  not g13287 (n_6737, n7191);
  and g13288 (n7192, n983, n_6737);
  not g13289 (n_6738, n7192);
  and g13290 (n7193, n987, n_6738);
  not g13291 (n_6739, n7193);
  and g13292 (n7194, n991, n_6739);
  not g13293 (n_6740, n7194);
  and g13294 (n7195, n995, n_6740);
  not g13295 (n_6741, n7195);
  and g13296 (n7196, n999, n_6741);
  not g13297 (n_6742, n7196);
  and g13298 (n7197, n1003, n_6742);
  not g13299 (n_6743, n7197);
  and g13300 (n7198, n1007, n_6743);
  not g13301 (n_6744, n7198);
  and g13302 (n7199, n1011, n_6744);
  not g13303 (n_6745, n7199);
  and g13304 (n7200, n1015, n_6745);
  not g13305 (n_6746, n7200);
  and g13306 (n7201, n1019, n_6746);
  not g13307 (n_6747, n7201);
  and g13308 (n7202, n1023, n_6747);
  not g13309 (n_6748, n7202);
  and g13310 (n7203, n1027, n_6748);
  not g13311 (n_6749, n7203);
  and g13312 (n7204, n1031, n_6749);
  not g13313 (n_6750, n7204);
  and g13314 (n7205, n1035, n_6750);
  not g13315 (n_6751, n7205);
  and g13316 (n7206, n1039, n_6751);
  not g13317 (n_6752, n7206);
  and g13318 (n7207, n1043, n_6752);
  not g13319 (n_6753, n7207);
  and g13320 (n7208, n1047, n_6753);
  not g13321 (n_6754, n7208);
  and g13322 (n7209, n1051, n_6754);
  not g13323 (n_6755, n7209);
  and g13324 (n7210, n1055, n_6755);
  not g13325 (n_6756, n7210);
  and g13326 (n7211, n1059, n_6756);
  not g13327 (n_6757, n7211);
  and g13328 (n7212, n1574, n_6757);
  not g13329 (n_6758, n7212);
  and g13330 (n7213, n1576, n_6758);
  not g13331 (n_6759, n7213);
  and g13332 (n7214, n1837, n_6759);
  not g13333 (n_6760, n7214);
  and g13334 (n7215, n1068, n_6760);
  not g13335 (n_6761, n7215);
  and g13336 (n7216, n1072, n_6761);
  not g13337 (n_6762, n7216);
  and g13338 (n7217, n1076, n_6762);
  not g13339 (n_6763, n7217);
  and g13340 (n7218, n1080, n_6763);
  not g13341 (n_6764, n7218);
  and g13342 (n7219, n1084, n_6764);
  not g13343 (n_6765, n7219);
  and g13344 (n7220, n1088, n_6765);
  not g13345 (n_6766, n7220);
  and g13346 (n7221, n1092, n_6766);
  not g13347 (n_6767, n7221);
  and g13348 (n7222, n1096, n_6767);
  not g13349 (n_6768, n7222);
  and g13350 (n7223, n1100, n_6768);
  not g13351 (n_6769, n7223);
  and g13352 (n7224, n1104, n_6769);
  not g13353 (n_6770, n7224);
  and g13354 (n7225, n1108, n_6770);
  not g13355 (n_6771, n7225);
  and g13356 (n7226, n1112, n_6771);
  not g13357 (n_6772, n7226);
  and g13358 (n7227, n1116, n_6772);
  not g13359 (n_6773, n7227);
  and g13360 (n7228, n1120, n_6773);
  not g13361 (n_6774, n7228);
  and g13362 (n7229, n1124, n_6774);
  not g13363 (n_6775, n7229);
  and g13364 (n7230, n1128, n_6775);
  not g13365 (n_6776, n7230);
  and g13366 (n7231, n1132, n_6776);
  not g13367 (n_6777, n7231);
  and g13368 (n7232, n1136, n_6777);
  not g13369 (n_6778, n7232);
  and g13370 (n7233, n1140, n_6778);
  not g13371 (n_6779, n7233);
  and g13372 (n7234, n1144, n_6779);
  not g13373 (n_6780, n7234);
  and g13374 (n7235, n1148, n_6780);
  not g13375 (n_6781, n7235);
  and g13376 (n7236, n1152, n_6781);
  not g13377 (n_6782, n7236);
  and g13378 (n7237, n1156, n_6782);
  not g13379 (n_6783, n7237);
  and g13380 (n7238, n1160, n_6783);
  not g13381 (n_6784, n7238);
  and g13382 (n7239, n1164, n_6784);
  not g13383 (n_6785, n7239);
  and g13384 (n7240, n1168, n_6785);
  not g13385 (n_6786, n7240);
  and g13386 (n7241, n1172, n_6786);
  not g13387 (n_6787, n7241);
  and g13388 (n7242, n1176, n_6787);
  not g13389 (n_6788, n7242);
  and g13390 (n7243, n1180, n_6788);
  not g13391 (n_6789, n7243);
  and g13392 (n7244, n1184, n_6789);
  not g13393 (n_6790, n7244);
  and g13394 (n7245, n1188, n_6790);
  not g13395 (n_6791, n7245);
  and g13396 (n7246, n1192, n_6791);
  not g13397 (n_6792, n7246);
  and g13398 (n7247, n1196, n_6792);
  not g13399 (n_6793, n7247);
  and g13400 (n7248, n1200, n_6793);
  not g13401 (n_6794, n7248);
  and g13402 (n7249, n1204, n_6794);
  not g13403 (n_6795, n7249);
  and g13404 (n7250, n1208, n_6795);
  not g13405 (n_6796, n7250);
  and g13406 (n7251, n1212, n_6796);
  not g13407 (n_6797, n7251);
  and g13408 (n7252, n1216, n_6797);
  not g13409 (n_6798, n7252);
  and g13410 (n7253, n1220, n_6798);
  not g13411 (n_6799, n7253);
  and g13412 (n7254, n1224, n_6799);
  not g13413 (n_6800, n7254);
  and g13414 (n7255, n1228, n_6800);
  not g13415 (n_6801, n7255);
  and g13416 (n7256, n1232, n_6801);
  not g13417 (n_6802, n7256);
  and g13418 (n7257, n1236, n_6802);
  and g13419 (n7258, \req[70] , n_939);
  not g13420 (n_6803, n7257);
  and g13421 (\grant[70] , n_6803, n7258);
  not g13422 (n_6804, n575);
  and g13423 (n7260, n_6804, n1247);
  not g13424 (n_6805, n7260);
  and g13425 (n7261, n1252, n_6805);
  not g13426 (n_6806, n7261);
  and g13427 (n7262, n1256, n_6806);
  not g13428 (n_6807, n7262);
  and g13429 (n7263, n1260, n_6807);
  not g13430 (n_6808, n7263);
  and g13431 (n7264, n1264, n_6808);
  not g13432 (n_6809, n7264);
  and g13433 (n7265, n1268, n_6809);
  not g13434 (n_6810, n7265);
  and g13435 (n7266, n1272, n_6810);
  not g13436 (n_6811, n7266);
  and g13437 (n7267, n1276, n_6811);
  not g13438 (n_6812, n7267);
  and g13439 (n7268, n1280, n_6812);
  not g13440 (n_6813, n7268);
  and g13441 (n7269, n1284, n_6813);
  not g13442 (n_6814, n7269);
  and g13443 (n7270, n1288, n_6814);
  not g13444 (n_6815, n7270);
  and g13445 (n7271, n1292, n_6815);
  not g13446 (n_6816, n7271);
  and g13447 (n7272, n1296, n_6816);
  not g13448 (n_6817, n7272);
  and g13449 (n7273, n1300, n_6817);
  not g13450 (n_6818, n7273);
  and g13451 (n7274, n1304, n_6818);
  not g13452 (n_6819, n7274);
  and g13453 (n7275, n1308, n_6819);
  not g13454 (n_6820, n7275);
  and g13455 (n7276, n1312, n_6820);
  not g13456 (n_6821, n7276);
  and g13457 (n7277, n1316, n_6821);
  not g13458 (n_6822, n7277);
  and g13459 (n7278, n1320, n_6822);
  not g13460 (n_6823, n7278);
  and g13461 (n7279, n1324, n_6823);
  not g13462 (n_6824, n7279);
  and g13463 (n7280, n1328, n_6824);
  not g13464 (n_6825, n7280);
  and g13465 (n7281, n1332, n_6825);
  not g13466 (n_6826, n7281);
  and g13467 (n7282, n1336, n_6826);
  not g13468 (n_6827, n7282);
  and g13469 (n7283, n1340, n_6827);
  not g13470 (n_6828, n7283);
  and g13471 (n7284, n1344, n_6828);
  not g13472 (n_6829, n7284);
  and g13473 (n7285, n1348, n_6829);
  not g13474 (n_6830, n7285);
  and g13475 (n7286, n1352, n_6830);
  not g13476 (n_6831, n7286);
  and g13477 (n7287, n1356, n_6831);
  not g13478 (n_6832, n7287);
  and g13479 (n7288, n1360, n_6832);
  not g13480 (n_6833, n7288);
  and g13481 (n7289, n1364, n_6833);
  not g13482 (n_6834, n7289);
  and g13483 (n7290, n1368, n_6834);
  not g13484 (n_6835, n7290);
  and g13485 (n7291, n1372, n_6835);
  not g13486 (n_6836, n7291);
  and g13487 (n7292, n1376, n_6836);
  not g13488 (n_6837, n7292);
  and g13489 (n7293, n1380, n_6837);
  not g13490 (n_6838, n7293);
  and g13491 (n7294, n1384, n_6838);
  not g13492 (n_6839, n7294);
  and g13493 (n7295, n1388, n_6839);
  not g13494 (n_6840, n7295);
  and g13495 (n7296, n1392, n_6840);
  not g13496 (n_6841, n7296);
  and g13497 (n7297, n1396, n_6841);
  not g13498 (n_6842, n7297);
  and g13499 (n7298, n1663, n_6842);
  not g13500 (n_6843, n7298);
  and g13501 (n7299, n392, n_6843);
  not g13502 (n_6844, n7299);
  and g13503 (n7300, n396, n_6844);
  not g13504 (n_6845, n7300);
  and g13505 (n7301, n400, n_6845);
  not g13506 (n_6846, n7301);
  and g13507 (n7302, n404, n_6846);
  not g13508 (n_6847, n7302);
  and g13509 (n7303, n408, n_6847);
  not g13510 (n_6848, n7303);
  and g13511 (n7304, n412, n_6848);
  not g13512 (n_6849, n7304);
  and g13513 (n7305, n416, n_6849);
  not g13514 (n_6850, n7305);
  and g13515 (n7306, n420, n_6850);
  not g13516 (n_6851, n7306);
  and g13517 (n7307, n424, n_6851);
  not g13518 (n_6852, n7307);
  and g13519 (n7308, n428, n_6852);
  not g13520 (n_6853, n7308);
  and g13521 (n7309, n432, n_6853);
  not g13522 (n_6854, n7309);
  and g13523 (n7310, n436, n_6854);
  not g13524 (n_6855, n7310);
  and g13525 (n7311, n440, n_6855);
  not g13526 (n_6856, n7311);
  and g13527 (n7312, n444, n_6856);
  not g13528 (n_6857, n7312);
  and g13529 (n7313, n448, n_6857);
  not g13530 (n_6858, n7313);
  and g13531 (n7314, n452, n_6858);
  not g13532 (n_6859, n7314);
  and g13533 (n7315, n456, n_6859);
  not g13534 (n_6860, n7315);
  and g13535 (n7316, n460, n_6860);
  not g13536 (n_6861, n7316);
  and g13537 (n7317, n464, n_6861);
  not g13538 (n_6862, n7317);
  and g13539 (n7318, n468, n_6862);
  not g13540 (n_6863, n7318);
  and g13541 (n7319, n472, n_6863);
  not g13542 (n_6864, n7319);
  and g13543 (n7320, n476, n_6864);
  not g13544 (n_6865, n7320);
  and g13545 (n7321, n480, n_6865);
  not g13546 (n_6866, n7321);
  and g13547 (n7322, n484, n_6866);
  not g13548 (n_6867, n7322);
  and g13549 (n7323, n488, n_6867);
  not g13550 (n_6868, n7323);
  and g13551 (n7324, n492, n_6868);
  not g13552 (n_6869, n7324);
  and g13553 (n7325, n496, n_6869);
  not g13554 (n_6870, n7325);
  and g13555 (n7326, n500, n_6870);
  not g13556 (n_6871, n7326);
  and g13557 (n7327, n504, n_6871);
  not g13558 (n_6872, n7327);
  and g13559 (n7328, n508, n_6872);
  not g13560 (n_6873, n7328);
  and g13561 (n7329, n512, n_6873);
  not g13562 (n_6874, n7329);
  and g13563 (n7330, n516, n_6874);
  not g13564 (n_6875, n7330);
  and g13565 (n7331, n520, n_6875);
  not g13566 (n_6876, n7331);
  and g13567 (n7332, n524, n_6876);
  not g13568 (n_6877, n7332);
  and g13569 (n7333, n528, n_6877);
  not g13570 (n_6878, n7333);
  and g13571 (n7334, n532, n_6878);
  not g13572 (n_6879, n7334);
  and g13573 (n7335, n536, n_6879);
  not g13574 (n_6880, n7335);
  and g13575 (n7336, n540, n_6880);
  not g13576 (n_6881, n7336);
  and g13577 (n7337, n544, n_6881);
  not g13578 (n_6882, n7337);
  and g13579 (n7338, n548, n_6882);
  not g13580 (n_6883, n7338);
  and g13581 (n7339, n552, n_6883);
  not g13582 (n_6884, n7339);
  and g13583 (n7340, n556, n_6884);
  not g13584 (n_6885, n7340);
  and g13585 (n7341, n560, n_6885);
  not g13586 (n_6886, n7341);
  and g13587 (n7342, n564, n_6886);
  not g13588 (n_6887, n7342);
  and g13589 (n7343, n568, n_6887);
  and g13590 (n7344, \req[71] , n_332);
  not g13591 (n_6888, n7343);
  and g13592 (\grant[71] , n_6888, n7344);
  not g13593 (n_6889, n914);
  and g13594 (n7346, n579, n_6889);
  not g13595 (n_6890, n7346);
  and g13596 (n7347, n584, n_6890);
  not g13597 (n_6891, n7347);
  and g13598 (n7348, n588, n_6891);
  not g13599 (n_6892, n7348);
  and g13600 (n7349, n592, n_6892);
  not g13601 (n_6893, n7349);
  and g13602 (n7350, n596, n_6893);
  not g13603 (n_6894, n7350);
  and g13604 (n7351, n600, n_6894);
  not g13605 (n_6895, n7351);
  and g13606 (n7352, n604, n_6895);
  not g13607 (n_6896, n7352);
  and g13608 (n7353, n608, n_6896);
  not g13609 (n_6897, n7353);
  and g13610 (n7354, n612, n_6897);
  not g13611 (n_6898, n7354);
  and g13612 (n7355, n616, n_6898);
  not g13613 (n_6899, n7355);
  and g13614 (n7356, n620, n_6899);
  not g13615 (n_6900, n7356);
  and g13616 (n7357, n624, n_6900);
  not g13617 (n_6901, n7357);
  and g13618 (n7358, n628, n_6901);
  not g13619 (n_6902, n7358);
  and g13620 (n7359, n632, n_6902);
  not g13621 (n_6903, n7359);
  and g13622 (n7360, n636, n_6903);
  not g13623 (n_6904, n7360);
  and g13624 (n7361, n640, n_6904);
  not g13625 (n_6905, n7361);
  and g13626 (n7362, n644, n_6905);
  not g13627 (n_6906, n7362);
  and g13628 (n7363, n648, n_6906);
  not g13629 (n_6907, n7363);
  and g13630 (n7364, n652, n_6907);
  not g13631 (n_6908, n7364);
  and g13632 (n7365, n656, n_6908);
  not g13633 (n_6909, n7365);
  and g13634 (n7366, n660, n_6909);
  not g13635 (n_6910, n7366);
  and g13636 (n7367, n664, n_6910);
  not g13637 (n_6911, n7367);
  and g13638 (n7368, n668, n_6911);
  not g13639 (n_6912, n7368);
  and g13640 (n7369, n672, n_6912);
  not g13641 (n_6913, n7369);
  and g13642 (n7370, n676, n_6913);
  not g13643 (n_6914, n7370);
  and g13644 (n7371, n680, n_6914);
  not g13645 (n_6915, n7371);
  and g13646 (n7372, n684, n_6915);
  not g13647 (n_6916, n7372);
  and g13648 (n7373, n688, n_6916);
  not g13649 (n_6917, n7373);
  and g13650 (n7374, n692, n_6917);
  not g13651 (n_6918, n7374);
  and g13652 (n7375, n696, n_6918);
  not g13653 (n_6919, n7375);
  and g13654 (n7376, n700, n_6919);
  not g13655 (n_6920, n7376);
  and g13656 (n7377, n704, n_6920);
  not g13657 (n_6921, n7377);
  and g13658 (n7378, n708, n_6921);
  not g13659 (n_6922, n7378);
  and g13660 (n7379, n712, n_6922);
  not g13661 (n_6923, n7379);
  and g13662 (n7380, n716, n_6923);
  not g13663 (n_6924, n7380);
  and g13664 (n7381, n720, n_6924);
  not g13665 (n_6925, n7381);
  and g13666 (n7382, n1484, n_6925);
  not g13667 (n_6926, n7382);
  and g13668 (n7383, n1486, n_6926);
  not g13669 (n_6927, n7383);
  and g13670 (n7384, n1750, n_6927);
  not g13671 (n_6928, n7384);
  and g13672 (n7385, n731, n_6928);
  not g13673 (n_6929, n7385);
  and g13674 (n7386, n735, n_6929);
  not g13675 (n_6930, n7386);
  and g13676 (n7387, n739, n_6930);
  not g13677 (n_6931, n7387);
  and g13678 (n7388, n743, n_6931);
  not g13679 (n_6932, n7388);
  and g13680 (n7389, n747, n_6932);
  not g13681 (n_6933, n7389);
  and g13682 (n7390, n751, n_6933);
  not g13683 (n_6934, n7390);
  and g13684 (n7391, n755, n_6934);
  not g13685 (n_6935, n7391);
  and g13686 (n7392, n759, n_6935);
  not g13687 (n_6936, n7392);
  and g13688 (n7393, n763, n_6936);
  not g13689 (n_6937, n7393);
  and g13690 (n7394, n767, n_6937);
  not g13691 (n_6938, n7394);
  and g13692 (n7395, n771, n_6938);
  not g13693 (n_6939, n7395);
  and g13694 (n7396, n775, n_6939);
  not g13695 (n_6940, n7396);
  and g13696 (n7397, n779, n_6940);
  not g13697 (n_6941, n7397);
  and g13698 (n7398, n783, n_6941);
  not g13699 (n_6942, n7398);
  and g13700 (n7399, n787, n_6942);
  not g13701 (n_6943, n7399);
  and g13702 (n7400, n791, n_6943);
  not g13703 (n_6944, n7400);
  and g13704 (n7401, n795, n_6944);
  not g13705 (n_6945, n7401);
  and g13706 (n7402, n799, n_6945);
  not g13707 (n_6946, n7402);
  and g13708 (n7403, n803, n_6946);
  not g13709 (n_6947, n7403);
  and g13710 (n7404, n807, n_6947);
  not g13711 (n_6948, n7404);
  and g13712 (n7405, n811, n_6948);
  not g13713 (n_6949, n7405);
  and g13714 (n7406, n815, n_6949);
  not g13715 (n_6950, n7406);
  and g13716 (n7407, n819, n_6950);
  not g13717 (n_6951, n7407);
  and g13718 (n7408, n823, n_6951);
  not g13719 (n_6952, n7408);
  and g13720 (n7409, n827, n_6952);
  not g13721 (n_6953, n7409);
  and g13722 (n7410, n831, n_6953);
  not g13723 (n_6954, n7410);
  and g13724 (n7411, n835, n_6954);
  not g13725 (n_6955, n7411);
  and g13726 (n7412, n839, n_6955);
  not g13727 (n_6956, n7412);
  and g13728 (n7413, n843, n_6956);
  not g13729 (n_6957, n7413);
  and g13730 (n7414, n847, n_6957);
  not g13731 (n_6958, n7414);
  and g13732 (n7415, n851, n_6958);
  not g13733 (n_6959, n7415);
  and g13734 (n7416, n855, n_6959);
  not g13735 (n_6960, n7416);
  and g13736 (n7417, n859, n_6960);
  not g13737 (n_6961, n7417);
  and g13738 (n7418, n863, n_6961);
  not g13739 (n_6962, n7418);
  and g13740 (n7419, n867, n_6962);
  not g13741 (n_6963, n7419);
  and g13742 (n7420, n871, n_6963);
  not g13743 (n_6964, n7420);
  and g13744 (n7421, n875, n_6964);
  not g13745 (n_6965, n7421);
  and g13746 (n7422, n879, n_6965);
  not g13747 (n_6966, n7422);
  and g13748 (n7423, n883, n_6966);
  not g13749 (n_6967, n7423);
  and g13750 (n7424, n887, n_6967);
  not g13751 (n_6968, n7424);
  and g13752 (n7425, n891, n_6968);
  not g13753 (n_6969, n7425);
  and g13754 (n7426, n895, n_6969);
  not g13755 (n_6970, n7426);
  and g13756 (n7427, n899, n_6970);
  not g13757 (n_6971, n7427);
  and g13758 (n7428, n903, n_6971);
  not g13759 (n_6972, n7428);
  and g13760 (n7429, n907, n_6972);
  and g13761 (n7430, \req[72] , n_737);
  not g13762 (n_6973, n7429);
  and g13763 (\grant[72] , n_6973, n7430);
  not g13764 (n_6974, n1251);
  and g13765 (n7432, n918, n_6974);
  not g13766 (n_6975, n7432);
  and g13767 (n7433, n923, n_6975);
  not g13768 (n_6976, n7433);
  and g13769 (n7434, n927, n_6976);
  not g13770 (n_6977, n7434);
  and g13771 (n7435, n931, n_6977);
  not g13772 (n_6978, n7435);
  and g13773 (n7436, n935, n_6978);
  not g13774 (n_6979, n7436);
  and g13775 (n7437, n939, n_6979);
  not g13776 (n_6980, n7437);
  and g13777 (n7438, n943, n_6980);
  not g13778 (n_6981, n7438);
  and g13779 (n7439, n947, n_6981);
  not g13780 (n_6982, n7439);
  and g13781 (n7440, n951, n_6982);
  not g13782 (n_6983, n7440);
  and g13783 (n7441, n955, n_6983);
  not g13784 (n_6984, n7441);
  and g13785 (n7442, n959, n_6984);
  not g13786 (n_6985, n7442);
  and g13787 (n7443, n963, n_6985);
  not g13788 (n_6986, n7443);
  and g13789 (n7444, n967, n_6986);
  not g13790 (n_6987, n7444);
  and g13791 (n7445, n971, n_6987);
  not g13792 (n_6988, n7445);
  and g13793 (n7446, n975, n_6988);
  not g13794 (n_6989, n7446);
  and g13795 (n7447, n979, n_6989);
  not g13796 (n_6990, n7447);
  and g13797 (n7448, n983, n_6990);
  not g13798 (n_6991, n7448);
  and g13799 (n7449, n987, n_6991);
  not g13800 (n_6992, n7449);
  and g13801 (n7450, n991, n_6992);
  not g13802 (n_6993, n7450);
  and g13803 (n7451, n995, n_6993);
  not g13804 (n_6994, n7451);
  and g13805 (n7452, n999, n_6994);
  not g13806 (n_6995, n7452);
  and g13807 (n7453, n1003, n_6995);
  not g13808 (n_6996, n7453);
  and g13809 (n7454, n1007, n_6996);
  not g13810 (n_6997, n7454);
  and g13811 (n7455, n1011, n_6997);
  not g13812 (n_6998, n7455);
  and g13813 (n7456, n1015, n_6998);
  not g13814 (n_6999, n7456);
  and g13815 (n7457, n1019, n_6999);
  not g13816 (n_7000, n7457);
  and g13817 (n7458, n1023, n_7000);
  not g13818 (n_7001, n7458);
  and g13819 (n7459, n1027, n_7001);
  not g13820 (n_7002, n7459);
  and g13821 (n7460, n1031, n_7002);
  not g13822 (n_7003, n7460);
  and g13823 (n7461, n1035, n_7003);
  not g13824 (n_7004, n7461);
  and g13825 (n7462, n1039, n_7004);
  not g13826 (n_7005, n7462);
  and g13827 (n7463, n1043, n_7005);
  not g13828 (n_7006, n7463);
  and g13829 (n7464, n1047, n_7006);
  not g13830 (n_7007, n7464);
  and g13831 (n7465, n1051, n_7007);
  not g13832 (n_7008, n7465);
  and g13833 (n7466, n1055, n_7008);
  not g13834 (n_7009, n7466);
  and g13835 (n7467, n1059, n_7009);
  not g13836 (n_7010, n7467);
  and g13837 (n7468, n1574, n_7010);
  not g13838 (n_7011, n7468);
  and g13839 (n7469, n1576, n_7011);
  not g13840 (n_7012, n7469);
  and g13841 (n7470, n1837, n_7012);
  not g13842 (n_7013, n7470);
  and g13843 (n7471, n1068, n_7013);
  not g13844 (n_7014, n7471);
  and g13845 (n7472, n1072, n_7014);
  not g13846 (n_7015, n7472);
  and g13847 (n7473, n1076, n_7015);
  not g13848 (n_7016, n7473);
  and g13849 (n7474, n1080, n_7016);
  not g13850 (n_7017, n7474);
  and g13851 (n7475, n1084, n_7017);
  not g13852 (n_7018, n7475);
  and g13853 (n7476, n1088, n_7018);
  not g13854 (n_7019, n7476);
  and g13855 (n7477, n1092, n_7019);
  not g13856 (n_7020, n7477);
  and g13857 (n7478, n1096, n_7020);
  not g13858 (n_7021, n7478);
  and g13859 (n7479, n1100, n_7021);
  not g13860 (n_7022, n7479);
  and g13861 (n7480, n1104, n_7022);
  not g13862 (n_7023, n7480);
  and g13863 (n7481, n1108, n_7023);
  not g13864 (n_7024, n7481);
  and g13865 (n7482, n1112, n_7024);
  not g13866 (n_7025, n7482);
  and g13867 (n7483, n1116, n_7025);
  not g13868 (n_7026, n7483);
  and g13869 (n7484, n1120, n_7026);
  not g13870 (n_7027, n7484);
  and g13871 (n7485, n1124, n_7027);
  not g13872 (n_7028, n7485);
  and g13873 (n7486, n1128, n_7028);
  not g13874 (n_7029, n7486);
  and g13875 (n7487, n1132, n_7029);
  not g13876 (n_7030, n7487);
  and g13877 (n7488, n1136, n_7030);
  not g13878 (n_7031, n7488);
  and g13879 (n7489, n1140, n_7031);
  not g13880 (n_7032, n7489);
  and g13881 (n7490, n1144, n_7032);
  not g13882 (n_7033, n7490);
  and g13883 (n7491, n1148, n_7033);
  not g13884 (n_7034, n7491);
  and g13885 (n7492, n1152, n_7034);
  not g13886 (n_7035, n7492);
  and g13887 (n7493, n1156, n_7035);
  not g13888 (n_7036, n7493);
  and g13889 (n7494, n1160, n_7036);
  not g13890 (n_7037, n7494);
  and g13891 (n7495, n1164, n_7037);
  not g13892 (n_7038, n7495);
  and g13893 (n7496, n1168, n_7038);
  not g13894 (n_7039, n7496);
  and g13895 (n7497, n1172, n_7039);
  not g13896 (n_7040, n7497);
  and g13897 (n7498, n1176, n_7040);
  not g13898 (n_7041, n7498);
  and g13899 (n7499, n1180, n_7041);
  not g13900 (n_7042, n7499);
  and g13901 (n7500, n1184, n_7042);
  not g13902 (n_7043, n7500);
  and g13903 (n7501, n1188, n_7043);
  not g13904 (n_7044, n7501);
  and g13905 (n7502, n1192, n_7044);
  not g13906 (n_7045, n7502);
  and g13907 (n7503, n1196, n_7045);
  not g13908 (n_7046, n7503);
  and g13909 (n7504, n1200, n_7046);
  not g13910 (n_7047, n7504);
  and g13911 (n7505, n1204, n_7047);
  not g13912 (n_7048, n7505);
  and g13913 (n7506, n1208, n_7048);
  not g13914 (n_7049, n7506);
  and g13915 (n7507, n1212, n_7049);
  not g13916 (n_7050, n7507);
  and g13917 (n7508, n1216, n_7050);
  not g13918 (n_7051, n7508);
  and g13919 (n7509, n1220, n_7051);
  not g13920 (n_7052, n7509);
  and g13921 (n7510, n1224, n_7052);
  not g13922 (n_7053, n7510);
  and g13923 (n7511, n1228, n_7053);
  not g13924 (n_7054, n7511);
  and g13925 (n7512, n1232, n_7054);
  not g13926 (n_7055, n7512);
  and g13927 (n7513, n1236, n_7055);
  not g13928 (n_7056, n7513);
  and g13929 (n7514, n1240, n_7056);
  not g13930 (n_7057, n7514);
  and g13931 (n7515, n1244, n_7057);
  and g13932 (n7516, \req[73] , n_943);
  not g13933 (n_7058, n7515);
  and g13934 (\grant[73] , n_7058, n7516);
  not g13935 (n_7059, n583);
  and g13936 (n7518, n_7059, n1255);
  not g13937 (n_7060, n7518);
  and g13938 (n7519, n1260, n_7060);
  not g13939 (n_7061, n7519);
  and g13940 (n7520, n1264, n_7061);
  not g13941 (n_7062, n7520);
  and g13942 (n7521, n1268, n_7062);
  not g13943 (n_7063, n7521);
  and g13944 (n7522, n1272, n_7063);
  not g13945 (n_7064, n7522);
  and g13946 (n7523, n1276, n_7064);
  not g13947 (n_7065, n7523);
  and g13948 (n7524, n1280, n_7065);
  not g13949 (n_7066, n7524);
  and g13950 (n7525, n1284, n_7066);
  not g13951 (n_7067, n7525);
  and g13952 (n7526, n1288, n_7067);
  not g13953 (n_7068, n7526);
  and g13954 (n7527, n1292, n_7068);
  not g13955 (n_7069, n7527);
  and g13956 (n7528, n1296, n_7069);
  not g13957 (n_7070, n7528);
  and g13958 (n7529, n1300, n_7070);
  not g13959 (n_7071, n7529);
  and g13960 (n7530, n1304, n_7071);
  not g13961 (n_7072, n7530);
  and g13962 (n7531, n1308, n_7072);
  not g13963 (n_7073, n7531);
  and g13964 (n7532, n1312, n_7073);
  not g13965 (n_7074, n7532);
  and g13966 (n7533, n1316, n_7074);
  not g13967 (n_7075, n7533);
  and g13968 (n7534, n1320, n_7075);
  not g13969 (n_7076, n7534);
  and g13970 (n7535, n1324, n_7076);
  not g13971 (n_7077, n7535);
  and g13972 (n7536, n1328, n_7077);
  not g13973 (n_7078, n7536);
  and g13974 (n7537, n1332, n_7078);
  not g13975 (n_7079, n7537);
  and g13976 (n7538, n1336, n_7079);
  not g13977 (n_7080, n7538);
  and g13978 (n7539, n1340, n_7080);
  not g13979 (n_7081, n7539);
  and g13980 (n7540, n1344, n_7081);
  not g13981 (n_7082, n7540);
  and g13982 (n7541, n1348, n_7082);
  not g13983 (n_7083, n7541);
  and g13984 (n7542, n1352, n_7083);
  not g13985 (n_7084, n7542);
  and g13986 (n7543, n1356, n_7084);
  not g13987 (n_7085, n7543);
  and g13988 (n7544, n1360, n_7085);
  not g13989 (n_7086, n7544);
  and g13990 (n7545, n1364, n_7086);
  not g13991 (n_7087, n7545);
  and g13992 (n7546, n1368, n_7087);
  not g13993 (n_7088, n7546);
  and g13994 (n7547, n1372, n_7088);
  not g13995 (n_7089, n7547);
  and g13996 (n7548, n1376, n_7089);
  not g13997 (n_7090, n7548);
  and g13998 (n7549, n1380, n_7090);
  not g13999 (n_7091, n7549);
  and g14000 (n7550, n1384, n_7091);
  not g14001 (n_7092, n7550);
  and g14002 (n7551, n1388, n_7092);
  not g14003 (n_7093, n7551);
  and g14004 (n7552, n1392, n_7093);
  not g14005 (n_7094, n7552);
  and g14006 (n7553, n1396, n_7094);
  not g14007 (n_7095, n7553);
  and g14008 (n7554, n1663, n_7095);
  not g14009 (n_7096, n7554);
  and g14010 (n7555, n392, n_7096);
  not g14011 (n_7097, n7555);
  and g14012 (n7556, n396, n_7097);
  not g14013 (n_7098, n7556);
  and g14014 (n7557, n400, n_7098);
  not g14015 (n_7099, n7557);
  and g14016 (n7558, n404, n_7099);
  not g14017 (n_7100, n7558);
  and g14018 (n7559, n408, n_7100);
  not g14019 (n_7101, n7559);
  and g14020 (n7560, n412, n_7101);
  not g14021 (n_7102, n7560);
  and g14022 (n7561, n416, n_7102);
  not g14023 (n_7103, n7561);
  and g14024 (n7562, n420, n_7103);
  not g14025 (n_7104, n7562);
  and g14026 (n7563, n424, n_7104);
  not g14027 (n_7105, n7563);
  and g14028 (n7564, n428, n_7105);
  not g14029 (n_7106, n7564);
  and g14030 (n7565, n432, n_7106);
  not g14031 (n_7107, n7565);
  and g14032 (n7566, n436, n_7107);
  not g14033 (n_7108, n7566);
  and g14034 (n7567, n440, n_7108);
  not g14035 (n_7109, n7567);
  and g14036 (n7568, n444, n_7109);
  not g14037 (n_7110, n7568);
  and g14038 (n7569, n448, n_7110);
  not g14039 (n_7111, n7569);
  and g14040 (n7570, n452, n_7111);
  not g14041 (n_7112, n7570);
  and g14042 (n7571, n456, n_7112);
  not g14043 (n_7113, n7571);
  and g14044 (n7572, n460, n_7113);
  not g14045 (n_7114, n7572);
  and g14046 (n7573, n464, n_7114);
  not g14047 (n_7115, n7573);
  and g14048 (n7574, n468, n_7115);
  not g14049 (n_7116, n7574);
  and g14050 (n7575, n472, n_7116);
  not g14051 (n_7117, n7575);
  and g14052 (n7576, n476, n_7117);
  not g14053 (n_7118, n7576);
  and g14054 (n7577, n480, n_7118);
  not g14055 (n_7119, n7577);
  and g14056 (n7578, n484, n_7119);
  not g14057 (n_7120, n7578);
  and g14058 (n7579, n488, n_7120);
  not g14059 (n_7121, n7579);
  and g14060 (n7580, n492, n_7121);
  not g14061 (n_7122, n7580);
  and g14062 (n7581, n496, n_7122);
  not g14063 (n_7123, n7581);
  and g14064 (n7582, n500, n_7123);
  not g14065 (n_7124, n7582);
  and g14066 (n7583, n504, n_7124);
  not g14067 (n_7125, n7583);
  and g14068 (n7584, n508, n_7125);
  not g14069 (n_7126, n7584);
  and g14070 (n7585, n512, n_7126);
  not g14071 (n_7127, n7585);
  and g14072 (n7586, n516, n_7127);
  not g14073 (n_7128, n7586);
  and g14074 (n7587, n520, n_7128);
  not g14075 (n_7129, n7587);
  and g14076 (n7588, n524, n_7129);
  not g14077 (n_7130, n7588);
  and g14078 (n7589, n528, n_7130);
  not g14079 (n_7131, n7589);
  and g14080 (n7590, n532, n_7131);
  not g14081 (n_7132, n7590);
  and g14082 (n7591, n536, n_7132);
  not g14083 (n_7133, n7591);
  and g14084 (n7592, n540, n_7133);
  not g14085 (n_7134, n7592);
  and g14086 (n7593, n544, n_7134);
  not g14087 (n_7135, n7593);
  and g14088 (n7594, n548, n_7135);
  not g14089 (n_7136, n7594);
  and g14090 (n7595, n552, n_7136);
  not g14091 (n_7137, n7595);
  and g14092 (n7596, n556, n_7137);
  not g14093 (n_7138, n7596);
  and g14094 (n7597, n560, n_7138);
  not g14095 (n_7139, n7597);
  and g14096 (n7598, n564, n_7139);
  not g14097 (n_7140, n7598);
  and g14098 (n7599, n568, n_7140);
  not g14099 (n_7141, n7599);
  and g14100 (n7600, n572, n_7141);
  not g14101 (n_7142, n7600);
  and g14102 (n7601, n576, n_7142);
  and g14103 (n7602, \req[74] , n_346);
  not g14104 (n_7143, n7601);
  and g14105 (\grant[74] , n_7143, n7602);
  not g14106 (n_7144, n922);
  and g14107 (n7604, n587, n_7144);
  not g14108 (n_7145, n7604);
  and g14109 (n7605, n592, n_7145);
  not g14110 (n_7146, n7605);
  and g14111 (n7606, n596, n_7146);
  not g14112 (n_7147, n7606);
  and g14113 (n7607, n600, n_7147);
  not g14114 (n_7148, n7607);
  and g14115 (n7608, n604, n_7148);
  not g14116 (n_7149, n7608);
  and g14117 (n7609, n608, n_7149);
  not g14118 (n_7150, n7609);
  and g14119 (n7610, n612, n_7150);
  not g14120 (n_7151, n7610);
  and g14121 (n7611, n616, n_7151);
  not g14122 (n_7152, n7611);
  and g14123 (n7612, n620, n_7152);
  not g14124 (n_7153, n7612);
  and g14125 (n7613, n624, n_7153);
  not g14126 (n_7154, n7613);
  and g14127 (n7614, n628, n_7154);
  not g14128 (n_7155, n7614);
  and g14129 (n7615, n632, n_7155);
  not g14130 (n_7156, n7615);
  and g14131 (n7616, n636, n_7156);
  not g14132 (n_7157, n7616);
  and g14133 (n7617, n640, n_7157);
  not g14134 (n_7158, n7617);
  and g14135 (n7618, n644, n_7158);
  not g14136 (n_7159, n7618);
  and g14137 (n7619, n648, n_7159);
  not g14138 (n_7160, n7619);
  and g14139 (n7620, n652, n_7160);
  not g14140 (n_7161, n7620);
  and g14141 (n7621, n656, n_7161);
  not g14142 (n_7162, n7621);
  and g14143 (n7622, n660, n_7162);
  not g14144 (n_7163, n7622);
  and g14145 (n7623, n664, n_7163);
  not g14146 (n_7164, n7623);
  and g14147 (n7624, n668, n_7164);
  not g14148 (n_7165, n7624);
  and g14149 (n7625, n672, n_7165);
  not g14150 (n_7166, n7625);
  and g14151 (n7626, n676, n_7166);
  not g14152 (n_7167, n7626);
  and g14153 (n7627, n680, n_7167);
  not g14154 (n_7168, n7627);
  and g14155 (n7628, n684, n_7168);
  not g14156 (n_7169, n7628);
  and g14157 (n7629, n688, n_7169);
  not g14158 (n_7170, n7629);
  and g14159 (n7630, n692, n_7170);
  not g14160 (n_7171, n7630);
  and g14161 (n7631, n696, n_7171);
  not g14162 (n_7172, n7631);
  and g14163 (n7632, n700, n_7172);
  not g14164 (n_7173, n7632);
  and g14165 (n7633, n704, n_7173);
  not g14166 (n_7174, n7633);
  and g14167 (n7634, n708, n_7174);
  not g14168 (n_7175, n7634);
  and g14169 (n7635, n712, n_7175);
  not g14170 (n_7176, n7635);
  and g14171 (n7636, n716, n_7176);
  not g14172 (n_7177, n7636);
  and g14173 (n7637, n720, n_7177);
  not g14174 (n_7178, n7637);
  and g14175 (n7638, n1484, n_7178);
  not g14176 (n_7179, n7638);
  and g14177 (n7639, n1486, n_7179);
  not g14178 (n_7180, n7639);
  and g14179 (n7640, n1750, n_7180);
  not g14180 (n_7181, n7640);
  and g14181 (n7641, n731, n_7181);
  not g14182 (n_7182, n7641);
  and g14183 (n7642, n735, n_7182);
  not g14184 (n_7183, n7642);
  and g14185 (n7643, n739, n_7183);
  not g14186 (n_7184, n7643);
  and g14187 (n7644, n743, n_7184);
  not g14188 (n_7185, n7644);
  and g14189 (n7645, n747, n_7185);
  not g14190 (n_7186, n7645);
  and g14191 (n7646, n751, n_7186);
  not g14192 (n_7187, n7646);
  and g14193 (n7647, n755, n_7187);
  not g14194 (n_7188, n7647);
  and g14195 (n7648, n759, n_7188);
  not g14196 (n_7189, n7648);
  and g14197 (n7649, n763, n_7189);
  not g14198 (n_7190, n7649);
  and g14199 (n7650, n767, n_7190);
  not g14200 (n_7191, n7650);
  and g14201 (n7651, n771, n_7191);
  not g14202 (n_7192, n7651);
  and g14203 (n7652, n775, n_7192);
  not g14204 (n_7193, n7652);
  and g14205 (n7653, n779, n_7193);
  not g14206 (n_7194, n7653);
  and g14207 (n7654, n783, n_7194);
  not g14208 (n_7195, n7654);
  and g14209 (n7655, n787, n_7195);
  not g14210 (n_7196, n7655);
  and g14211 (n7656, n791, n_7196);
  not g14212 (n_7197, n7656);
  and g14213 (n7657, n795, n_7197);
  not g14214 (n_7198, n7657);
  and g14215 (n7658, n799, n_7198);
  not g14216 (n_7199, n7658);
  and g14217 (n7659, n803, n_7199);
  not g14218 (n_7200, n7659);
  and g14219 (n7660, n807, n_7200);
  not g14220 (n_7201, n7660);
  and g14221 (n7661, n811, n_7201);
  not g14222 (n_7202, n7661);
  and g14223 (n7662, n815, n_7202);
  not g14224 (n_7203, n7662);
  and g14225 (n7663, n819, n_7203);
  not g14226 (n_7204, n7663);
  and g14227 (n7664, n823, n_7204);
  not g14228 (n_7205, n7664);
  and g14229 (n7665, n827, n_7205);
  not g14230 (n_7206, n7665);
  and g14231 (n7666, n831, n_7206);
  not g14232 (n_7207, n7666);
  and g14233 (n7667, n835, n_7207);
  not g14234 (n_7208, n7667);
  and g14235 (n7668, n839, n_7208);
  not g14236 (n_7209, n7668);
  and g14237 (n7669, n843, n_7209);
  not g14238 (n_7210, n7669);
  and g14239 (n7670, n847, n_7210);
  not g14240 (n_7211, n7670);
  and g14241 (n7671, n851, n_7211);
  not g14242 (n_7212, n7671);
  and g14243 (n7672, n855, n_7212);
  not g14244 (n_7213, n7672);
  and g14245 (n7673, n859, n_7213);
  not g14246 (n_7214, n7673);
  and g14247 (n7674, n863, n_7214);
  not g14248 (n_7215, n7674);
  and g14249 (n7675, n867, n_7215);
  not g14250 (n_7216, n7675);
  and g14251 (n7676, n871, n_7216);
  not g14252 (n_7217, n7676);
  and g14253 (n7677, n875, n_7217);
  not g14254 (n_7218, n7677);
  and g14255 (n7678, n879, n_7218);
  not g14256 (n_7219, n7678);
  and g14257 (n7679, n883, n_7219);
  not g14258 (n_7220, n7679);
  and g14259 (n7680, n887, n_7220);
  not g14260 (n_7221, n7680);
  and g14261 (n7681, n891, n_7221);
  not g14262 (n_7222, n7681);
  and g14263 (n7682, n895, n_7222);
  not g14264 (n_7223, n7682);
  and g14265 (n7683, n899, n_7223);
  not g14266 (n_7224, n7683);
  and g14267 (n7684, n903, n_7224);
  not g14268 (n_7225, n7684);
  and g14269 (n7685, n907, n_7225);
  not g14270 (n_7226, n7685);
  and g14271 (n7686, n911, n_7226);
  not g14272 (n_7227, n7686);
  and g14273 (n7687, n915, n_7227);
  and g14274 (n7688, \req[75] , n_743);
  not g14275 (n_7228, n7687);
  and g14276 (\grant[75] , n_7228, n7688);
  not g14277 (n_7229, n1259);
  and g14278 (n7690, n926, n_7229);
  not g14279 (n_7230, n7690);
  and g14280 (n7691, n931, n_7230);
  not g14281 (n_7231, n7691);
  and g14282 (n7692, n935, n_7231);
  not g14283 (n_7232, n7692);
  and g14284 (n7693, n939, n_7232);
  not g14285 (n_7233, n7693);
  and g14286 (n7694, n943, n_7233);
  not g14287 (n_7234, n7694);
  and g14288 (n7695, n947, n_7234);
  not g14289 (n_7235, n7695);
  and g14290 (n7696, n951, n_7235);
  not g14291 (n_7236, n7696);
  and g14292 (n7697, n955, n_7236);
  not g14293 (n_7237, n7697);
  and g14294 (n7698, n959, n_7237);
  not g14295 (n_7238, n7698);
  and g14296 (n7699, n963, n_7238);
  not g14297 (n_7239, n7699);
  and g14298 (n7700, n967, n_7239);
  not g14299 (n_7240, n7700);
  and g14300 (n7701, n971, n_7240);
  not g14301 (n_7241, n7701);
  and g14302 (n7702, n975, n_7241);
  not g14303 (n_7242, n7702);
  and g14304 (n7703, n979, n_7242);
  not g14305 (n_7243, n7703);
  and g14306 (n7704, n983, n_7243);
  not g14307 (n_7244, n7704);
  and g14308 (n7705, n987, n_7244);
  not g14309 (n_7245, n7705);
  and g14310 (n7706, n991, n_7245);
  not g14311 (n_7246, n7706);
  and g14312 (n7707, n995, n_7246);
  not g14313 (n_7247, n7707);
  and g14314 (n7708, n999, n_7247);
  not g14315 (n_7248, n7708);
  and g14316 (n7709, n1003, n_7248);
  not g14317 (n_7249, n7709);
  and g14318 (n7710, n1007, n_7249);
  not g14319 (n_7250, n7710);
  and g14320 (n7711, n1011, n_7250);
  not g14321 (n_7251, n7711);
  and g14322 (n7712, n1015, n_7251);
  not g14323 (n_7252, n7712);
  and g14324 (n7713, n1019, n_7252);
  not g14325 (n_7253, n7713);
  and g14326 (n7714, n1023, n_7253);
  not g14327 (n_7254, n7714);
  and g14328 (n7715, n1027, n_7254);
  not g14329 (n_7255, n7715);
  and g14330 (n7716, n1031, n_7255);
  not g14331 (n_7256, n7716);
  and g14332 (n7717, n1035, n_7256);
  not g14333 (n_7257, n7717);
  and g14334 (n7718, n1039, n_7257);
  not g14335 (n_7258, n7718);
  and g14336 (n7719, n1043, n_7258);
  not g14337 (n_7259, n7719);
  and g14338 (n7720, n1047, n_7259);
  not g14339 (n_7260, n7720);
  and g14340 (n7721, n1051, n_7260);
  not g14341 (n_7261, n7721);
  and g14342 (n7722, n1055, n_7261);
  not g14343 (n_7262, n7722);
  and g14344 (n7723, n1059, n_7262);
  not g14345 (n_7263, n7723);
  and g14346 (n7724, n1574, n_7263);
  not g14347 (n_7264, n7724);
  and g14348 (n7725, n1576, n_7264);
  not g14349 (n_7265, n7725);
  and g14350 (n7726, n1837, n_7265);
  not g14351 (n_7266, n7726);
  and g14352 (n7727, n1068, n_7266);
  not g14353 (n_7267, n7727);
  and g14354 (n7728, n1072, n_7267);
  not g14355 (n_7268, n7728);
  and g14356 (n7729, n1076, n_7268);
  not g14357 (n_7269, n7729);
  and g14358 (n7730, n1080, n_7269);
  not g14359 (n_7270, n7730);
  and g14360 (n7731, n1084, n_7270);
  not g14361 (n_7271, n7731);
  and g14362 (n7732, n1088, n_7271);
  not g14363 (n_7272, n7732);
  and g14364 (n7733, n1092, n_7272);
  not g14365 (n_7273, n7733);
  and g14366 (n7734, n1096, n_7273);
  not g14367 (n_7274, n7734);
  and g14368 (n7735, n1100, n_7274);
  not g14369 (n_7275, n7735);
  and g14370 (n7736, n1104, n_7275);
  not g14371 (n_7276, n7736);
  and g14372 (n7737, n1108, n_7276);
  not g14373 (n_7277, n7737);
  and g14374 (n7738, n1112, n_7277);
  not g14375 (n_7278, n7738);
  and g14376 (n7739, n1116, n_7278);
  not g14377 (n_7279, n7739);
  and g14378 (n7740, n1120, n_7279);
  not g14379 (n_7280, n7740);
  and g14380 (n7741, n1124, n_7280);
  not g14381 (n_7281, n7741);
  and g14382 (n7742, n1128, n_7281);
  not g14383 (n_7282, n7742);
  and g14384 (n7743, n1132, n_7282);
  not g14385 (n_7283, n7743);
  and g14386 (n7744, n1136, n_7283);
  not g14387 (n_7284, n7744);
  and g14388 (n7745, n1140, n_7284);
  not g14389 (n_7285, n7745);
  and g14390 (n7746, n1144, n_7285);
  not g14391 (n_7286, n7746);
  and g14392 (n7747, n1148, n_7286);
  not g14393 (n_7287, n7747);
  and g14394 (n7748, n1152, n_7287);
  not g14395 (n_7288, n7748);
  and g14396 (n7749, n1156, n_7288);
  not g14397 (n_7289, n7749);
  and g14398 (n7750, n1160, n_7289);
  not g14399 (n_7290, n7750);
  and g14400 (n7751, n1164, n_7290);
  not g14401 (n_7291, n7751);
  and g14402 (n7752, n1168, n_7291);
  not g14403 (n_7292, n7752);
  and g14404 (n7753, n1172, n_7292);
  not g14405 (n_7293, n7753);
  and g14406 (n7754, n1176, n_7293);
  not g14407 (n_7294, n7754);
  and g14408 (n7755, n1180, n_7294);
  not g14409 (n_7295, n7755);
  and g14410 (n7756, n1184, n_7295);
  not g14411 (n_7296, n7756);
  and g14412 (n7757, n1188, n_7296);
  not g14413 (n_7297, n7757);
  and g14414 (n7758, n1192, n_7297);
  not g14415 (n_7298, n7758);
  and g14416 (n7759, n1196, n_7298);
  not g14417 (n_7299, n7759);
  and g14418 (n7760, n1200, n_7299);
  not g14419 (n_7300, n7760);
  and g14420 (n7761, n1204, n_7300);
  not g14421 (n_7301, n7761);
  and g14422 (n7762, n1208, n_7301);
  not g14423 (n_7302, n7762);
  and g14424 (n7763, n1212, n_7302);
  not g14425 (n_7303, n7763);
  and g14426 (n7764, n1216, n_7303);
  not g14427 (n_7304, n7764);
  and g14428 (n7765, n1220, n_7304);
  not g14429 (n_7305, n7765);
  and g14430 (n7766, n1224, n_7305);
  not g14431 (n_7306, n7766);
  and g14432 (n7767, n1228, n_7306);
  not g14433 (n_7307, n7767);
  and g14434 (n7768, n1232, n_7307);
  not g14435 (n_7308, n7768);
  and g14436 (n7769, n1236, n_7308);
  not g14437 (n_7309, n7769);
  and g14438 (n7770, n1240, n_7309);
  not g14439 (n_7310, n7770);
  and g14440 (n7771, n1244, n_7310);
  not g14441 (n_7311, n7771);
  and g14442 (n7772, n1248, n_7311);
  not g14443 (n_7312, n7772);
  and g14444 (n7773, n1252, n_7312);
  and g14445 (n7774, \req[76] , n_947);
  not g14446 (n_7313, n7773);
  and g14447 (\grant[76] , n_7313, n7774);
  not g14448 (n_7314, n591);
  and g14449 (n7776, n_7314, n1263);
  not g14450 (n_7315, n7776);
  and g14451 (n7777, n1268, n_7315);
  not g14452 (n_7316, n7777);
  and g14453 (n7778, n1272, n_7316);
  not g14454 (n_7317, n7778);
  and g14455 (n7779, n1276, n_7317);
  not g14456 (n_7318, n7779);
  and g14457 (n7780, n1280, n_7318);
  not g14458 (n_7319, n7780);
  and g14459 (n7781, n1284, n_7319);
  not g14460 (n_7320, n7781);
  and g14461 (n7782, n1288, n_7320);
  not g14462 (n_7321, n7782);
  and g14463 (n7783, n1292, n_7321);
  not g14464 (n_7322, n7783);
  and g14465 (n7784, n1296, n_7322);
  not g14466 (n_7323, n7784);
  and g14467 (n7785, n1300, n_7323);
  not g14468 (n_7324, n7785);
  and g14469 (n7786, n1304, n_7324);
  not g14470 (n_7325, n7786);
  and g14471 (n7787, n1308, n_7325);
  not g14472 (n_7326, n7787);
  and g14473 (n7788, n1312, n_7326);
  not g14474 (n_7327, n7788);
  and g14475 (n7789, n1316, n_7327);
  not g14476 (n_7328, n7789);
  and g14477 (n7790, n1320, n_7328);
  not g14478 (n_7329, n7790);
  and g14479 (n7791, n1324, n_7329);
  not g14480 (n_7330, n7791);
  and g14481 (n7792, n1328, n_7330);
  not g14482 (n_7331, n7792);
  and g14483 (n7793, n1332, n_7331);
  not g14484 (n_7332, n7793);
  and g14485 (n7794, n1336, n_7332);
  not g14486 (n_7333, n7794);
  and g14487 (n7795, n1340, n_7333);
  not g14488 (n_7334, n7795);
  and g14489 (n7796, n1344, n_7334);
  not g14490 (n_7335, n7796);
  and g14491 (n7797, n1348, n_7335);
  not g14492 (n_7336, n7797);
  and g14493 (n7798, n1352, n_7336);
  not g14494 (n_7337, n7798);
  and g14495 (n7799, n1356, n_7337);
  not g14496 (n_7338, n7799);
  and g14497 (n7800, n1360, n_7338);
  not g14498 (n_7339, n7800);
  and g14499 (n7801, n1364, n_7339);
  not g14500 (n_7340, n7801);
  and g14501 (n7802, n1368, n_7340);
  not g14502 (n_7341, n7802);
  and g14503 (n7803, n1372, n_7341);
  not g14504 (n_7342, n7803);
  and g14505 (n7804, n1376, n_7342);
  not g14506 (n_7343, n7804);
  and g14507 (n7805, n1380, n_7343);
  not g14508 (n_7344, n7805);
  and g14509 (n7806, n1384, n_7344);
  not g14510 (n_7345, n7806);
  and g14511 (n7807, n1388, n_7345);
  not g14512 (n_7346, n7807);
  and g14513 (n7808, n1392, n_7346);
  not g14514 (n_7347, n7808);
  and g14515 (n7809, n1396, n_7347);
  not g14516 (n_7348, n7809);
  and g14517 (n7810, n1663, n_7348);
  not g14518 (n_7349, n7810);
  and g14519 (n7811, n392, n_7349);
  not g14520 (n_7350, n7811);
  and g14521 (n7812, n396, n_7350);
  not g14522 (n_7351, n7812);
  and g14523 (n7813, n400, n_7351);
  not g14524 (n_7352, n7813);
  and g14525 (n7814, n404, n_7352);
  not g14526 (n_7353, n7814);
  and g14527 (n7815, n408, n_7353);
  not g14528 (n_7354, n7815);
  and g14529 (n7816, n412, n_7354);
  not g14530 (n_7355, n7816);
  and g14531 (n7817, n416, n_7355);
  not g14532 (n_7356, n7817);
  and g14533 (n7818, n420, n_7356);
  not g14534 (n_7357, n7818);
  and g14535 (n7819, n424, n_7357);
  not g14536 (n_7358, n7819);
  and g14537 (n7820, n428, n_7358);
  not g14538 (n_7359, n7820);
  and g14539 (n7821, n432, n_7359);
  not g14540 (n_7360, n7821);
  and g14541 (n7822, n436, n_7360);
  not g14542 (n_7361, n7822);
  and g14543 (n7823, n440, n_7361);
  not g14544 (n_7362, n7823);
  and g14545 (n7824, n444, n_7362);
  not g14546 (n_7363, n7824);
  and g14547 (n7825, n448, n_7363);
  not g14548 (n_7364, n7825);
  and g14549 (n7826, n452, n_7364);
  not g14550 (n_7365, n7826);
  and g14551 (n7827, n456, n_7365);
  not g14552 (n_7366, n7827);
  and g14553 (n7828, n460, n_7366);
  not g14554 (n_7367, n7828);
  and g14555 (n7829, n464, n_7367);
  not g14556 (n_7368, n7829);
  and g14557 (n7830, n468, n_7368);
  not g14558 (n_7369, n7830);
  and g14559 (n7831, n472, n_7369);
  not g14560 (n_7370, n7831);
  and g14561 (n7832, n476, n_7370);
  not g14562 (n_7371, n7832);
  and g14563 (n7833, n480, n_7371);
  not g14564 (n_7372, n7833);
  and g14565 (n7834, n484, n_7372);
  not g14566 (n_7373, n7834);
  and g14567 (n7835, n488, n_7373);
  not g14568 (n_7374, n7835);
  and g14569 (n7836, n492, n_7374);
  not g14570 (n_7375, n7836);
  and g14571 (n7837, n496, n_7375);
  not g14572 (n_7376, n7837);
  and g14573 (n7838, n500, n_7376);
  not g14574 (n_7377, n7838);
  and g14575 (n7839, n504, n_7377);
  not g14576 (n_7378, n7839);
  and g14577 (n7840, n508, n_7378);
  not g14578 (n_7379, n7840);
  and g14579 (n7841, n512, n_7379);
  not g14580 (n_7380, n7841);
  and g14581 (n7842, n516, n_7380);
  not g14582 (n_7381, n7842);
  and g14583 (n7843, n520, n_7381);
  not g14584 (n_7382, n7843);
  and g14585 (n7844, n524, n_7382);
  not g14586 (n_7383, n7844);
  and g14587 (n7845, n528, n_7383);
  not g14588 (n_7384, n7845);
  and g14589 (n7846, n532, n_7384);
  not g14590 (n_7385, n7846);
  and g14591 (n7847, n536, n_7385);
  not g14592 (n_7386, n7847);
  and g14593 (n7848, n540, n_7386);
  not g14594 (n_7387, n7848);
  and g14595 (n7849, n544, n_7387);
  not g14596 (n_7388, n7849);
  and g14597 (n7850, n548, n_7388);
  not g14598 (n_7389, n7850);
  and g14599 (n7851, n552, n_7389);
  not g14600 (n_7390, n7851);
  and g14601 (n7852, n556, n_7390);
  not g14602 (n_7391, n7852);
  and g14603 (n7853, n560, n_7391);
  not g14604 (n_7392, n7853);
  and g14605 (n7854, n564, n_7392);
  not g14606 (n_7393, n7854);
  and g14607 (n7855, n568, n_7393);
  not g14608 (n_7394, n7855);
  and g14609 (n7856, n572, n_7394);
  not g14610 (n_7395, n7856);
  and g14611 (n7857, n576, n_7395);
  not g14612 (n_7396, n7857);
  and g14613 (n7858, n580, n_7396);
  not g14614 (n_7397, n7858);
  and g14615 (n7859, n584, n_7397);
  and g14616 (n7860, \req[77] , n_360);
  not g14617 (n_7398, n7859);
  and g14618 (\grant[77] , n_7398, n7860);
  not g14619 (n_7399, n930);
  and g14620 (n7862, n595, n_7399);
  not g14621 (n_7400, n7862);
  and g14622 (n7863, n600, n_7400);
  not g14623 (n_7401, n7863);
  and g14624 (n7864, n604, n_7401);
  not g14625 (n_7402, n7864);
  and g14626 (n7865, n608, n_7402);
  not g14627 (n_7403, n7865);
  and g14628 (n7866, n612, n_7403);
  not g14629 (n_7404, n7866);
  and g14630 (n7867, n616, n_7404);
  not g14631 (n_7405, n7867);
  and g14632 (n7868, n620, n_7405);
  not g14633 (n_7406, n7868);
  and g14634 (n7869, n624, n_7406);
  not g14635 (n_7407, n7869);
  and g14636 (n7870, n628, n_7407);
  not g14637 (n_7408, n7870);
  and g14638 (n7871, n632, n_7408);
  not g14639 (n_7409, n7871);
  and g14640 (n7872, n636, n_7409);
  not g14641 (n_7410, n7872);
  and g14642 (n7873, n640, n_7410);
  not g14643 (n_7411, n7873);
  and g14644 (n7874, n644, n_7411);
  not g14645 (n_7412, n7874);
  and g14646 (n7875, n648, n_7412);
  not g14647 (n_7413, n7875);
  and g14648 (n7876, n652, n_7413);
  not g14649 (n_7414, n7876);
  and g14650 (n7877, n656, n_7414);
  not g14651 (n_7415, n7877);
  and g14652 (n7878, n660, n_7415);
  not g14653 (n_7416, n7878);
  and g14654 (n7879, n664, n_7416);
  not g14655 (n_7417, n7879);
  and g14656 (n7880, n668, n_7417);
  not g14657 (n_7418, n7880);
  and g14658 (n7881, n672, n_7418);
  not g14659 (n_7419, n7881);
  and g14660 (n7882, n676, n_7419);
  not g14661 (n_7420, n7882);
  and g14662 (n7883, n680, n_7420);
  not g14663 (n_7421, n7883);
  and g14664 (n7884, n684, n_7421);
  not g14665 (n_7422, n7884);
  and g14666 (n7885, n688, n_7422);
  not g14667 (n_7423, n7885);
  and g14668 (n7886, n692, n_7423);
  not g14669 (n_7424, n7886);
  and g14670 (n7887, n696, n_7424);
  not g14671 (n_7425, n7887);
  and g14672 (n7888, n700, n_7425);
  not g14673 (n_7426, n7888);
  and g14674 (n7889, n704, n_7426);
  not g14675 (n_7427, n7889);
  and g14676 (n7890, n708, n_7427);
  not g14677 (n_7428, n7890);
  and g14678 (n7891, n712, n_7428);
  not g14679 (n_7429, n7891);
  and g14680 (n7892, n716, n_7429);
  not g14681 (n_7430, n7892);
  and g14682 (n7893, n720, n_7430);
  not g14683 (n_7431, n7893);
  and g14684 (n7894, n1484, n_7431);
  not g14685 (n_7432, n7894);
  and g14686 (n7895, n1486, n_7432);
  not g14687 (n_7433, n7895);
  and g14688 (n7896, n1750, n_7433);
  not g14689 (n_7434, n7896);
  and g14690 (n7897, n731, n_7434);
  not g14691 (n_7435, n7897);
  and g14692 (n7898, n735, n_7435);
  not g14693 (n_7436, n7898);
  and g14694 (n7899, n739, n_7436);
  not g14695 (n_7437, n7899);
  and g14696 (n7900, n743, n_7437);
  not g14697 (n_7438, n7900);
  and g14698 (n7901, n747, n_7438);
  not g14699 (n_7439, n7901);
  and g14700 (n7902, n751, n_7439);
  not g14701 (n_7440, n7902);
  and g14702 (n7903, n755, n_7440);
  not g14703 (n_7441, n7903);
  and g14704 (n7904, n759, n_7441);
  not g14705 (n_7442, n7904);
  and g14706 (n7905, n763, n_7442);
  not g14707 (n_7443, n7905);
  and g14708 (n7906, n767, n_7443);
  not g14709 (n_7444, n7906);
  and g14710 (n7907, n771, n_7444);
  not g14711 (n_7445, n7907);
  and g14712 (n7908, n775, n_7445);
  not g14713 (n_7446, n7908);
  and g14714 (n7909, n779, n_7446);
  not g14715 (n_7447, n7909);
  and g14716 (n7910, n783, n_7447);
  not g14717 (n_7448, n7910);
  and g14718 (n7911, n787, n_7448);
  not g14719 (n_7449, n7911);
  and g14720 (n7912, n791, n_7449);
  not g14721 (n_7450, n7912);
  and g14722 (n7913, n795, n_7450);
  not g14723 (n_7451, n7913);
  and g14724 (n7914, n799, n_7451);
  not g14725 (n_7452, n7914);
  and g14726 (n7915, n803, n_7452);
  not g14727 (n_7453, n7915);
  and g14728 (n7916, n807, n_7453);
  not g14729 (n_7454, n7916);
  and g14730 (n7917, n811, n_7454);
  not g14731 (n_7455, n7917);
  and g14732 (n7918, n815, n_7455);
  not g14733 (n_7456, n7918);
  and g14734 (n7919, n819, n_7456);
  not g14735 (n_7457, n7919);
  and g14736 (n7920, n823, n_7457);
  not g14737 (n_7458, n7920);
  and g14738 (n7921, n827, n_7458);
  not g14739 (n_7459, n7921);
  and g14740 (n7922, n831, n_7459);
  not g14741 (n_7460, n7922);
  and g14742 (n7923, n835, n_7460);
  not g14743 (n_7461, n7923);
  and g14744 (n7924, n839, n_7461);
  not g14745 (n_7462, n7924);
  and g14746 (n7925, n843, n_7462);
  not g14747 (n_7463, n7925);
  and g14748 (n7926, n847, n_7463);
  not g14749 (n_7464, n7926);
  and g14750 (n7927, n851, n_7464);
  not g14751 (n_7465, n7927);
  and g14752 (n7928, n855, n_7465);
  not g14753 (n_7466, n7928);
  and g14754 (n7929, n859, n_7466);
  not g14755 (n_7467, n7929);
  and g14756 (n7930, n863, n_7467);
  not g14757 (n_7468, n7930);
  and g14758 (n7931, n867, n_7468);
  not g14759 (n_7469, n7931);
  and g14760 (n7932, n871, n_7469);
  not g14761 (n_7470, n7932);
  and g14762 (n7933, n875, n_7470);
  not g14763 (n_7471, n7933);
  and g14764 (n7934, n879, n_7471);
  not g14765 (n_7472, n7934);
  and g14766 (n7935, n883, n_7472);
  not g14767 (n_7473, n7935);
  and g14768 (n7936, n887, n_7473);
  not g14769 (n_7474, n7936);
  and g14770 (n7937, n891, n_7474);
  not g14771 (n_7475, n7937);
  and g14772 (n7938, n895, n_7475);
  not g14773 (n_7476, n7938);
  and g14774 (n7939, n899, n_7476);
  not g14775 (n_7477, n7939);
  and g14776 (n7940, n903, n_7477);
  not g14777 (n_7478, n7940);
  and g14778 (n7941, n907, n_7478);
  not g14779 (n_7479, n7941);
  and g14780 (n7942, n911, n_7479);
  not g14781 (n_7480, n7942);
  and g14782 (n7943, n915, n_7480);
  not g14783 (n_7481, n7943);
  and g14784 (n7944, n919, n_7481);
  not g14785 (n_7482, n7944);
  and g14786 (n7945, n923, n_7482);
  and g14787 (n7946, \req[78] , n_749);
  not g14788 (n_7483, n7945);
  and g14789 (\grant[78] , n_7483, n7946);
  not g14790 (n_7484, n1267);
  and g14791 (n7948, n934, n_7484);
  not g14792 (n_7485, n7948);
  and g14793 (n7949, n939, n_7485);
  not g14794 (n_7486, n7949);
  and g14795 (n7950, n943, n_7486);
  not g14796 (n_7487, n7950);
  and g14797 (n7951, n947, n_7487);
  not g14798 (n_7488, n7951);
  and g14799 (n7952, n951, n_7488);
  not g14800 (n_7489, n7952);
  and g14801 (n7953, n955, n_7489);
  not g14802 (n_7490, n7953);
  and g14803 (n7954, n959, n_7490);
  not g14804 (n_7491, n7954);
  and g14805 (n7955, n963, n_7491);
  not g14806 (n_7492, n7955);
  and g14807 (n7956, n967, n_7492);
  not g14808 (n_7493, n7956);
  and g14809 (n7957, n971, n_7493);
  not g14810 (n_7494, n7957);
  and g14811 (n7958, n975, n_7494);
  not g14812 (n_7495, n7958);
  and g14813 (n7959, n979, n_7495);
  not g14814 (n_7496, n7959);
  and g14815 (n7960, n983, n_7496);
  not g14816 (n_7497, n7960);
  and g14817 (n7961, n987, n_7497);
  not g14818 (n_7498, n7961);
  and g14819 (n7962, n991, n_7498);
  not g14820 (n_7499, n7962);
  and g14821 (n7963, n995, n_7499);
  not g14822 (n_7500, n7963);
  and g14823 (n7964, n999, n_7500);
  not g14824 (n_7501, n7964);
  and g14825 (n7965, n1003, n_7501);
  not g14826 (n_7502, n7965);
  and g14827 (n7966, n1007, n_7502);
  not g14828 (n_7503, n7966);
  and g14829 (n7967, n1011, n_7503);
  not g14830 (n_7504, n7967);
  and g14831 (n7968, n1015, n_7504);
  not g14832 (n_7505, n7968);
  and g14833 (n7969, n1019, n_7505);
  not g14834 (n_7506, n7969);
  and g14835 (n7970, n1023, n_7506);
  not g14836 (n_7507, n7970);
  and g14837 (n7971, n1027, n_7507);
  not g14838 (n_7508, n7971);
  and g14839 (n7972, n1031, n_7508);
  not g14840 (n_7509, n7972);
  and g14841 (n7973, n1035, n_7509);
  not g14842 (n_7510, n7973);
  and g14843 (n7974, n1039, n_7510);
  not g14844 (n_7511, n7974);
  and g14845 (n7975, n1043, n_7511);
  not g14846 (n_7512, n7975);
  and g14847 (n7976, n1047, n_7512);
  not g14848 (n_7513, n7976);
  and g14849 (n7977, n1051, n_7513);
  not g14850 (n_7514, n7977);
  and g14851 (n7978, n1055, n_7514);
  not g14852 (n_7515, n7978);
  and g14853 (n7979, n1059, n_7515);
  not g14854 (n_7516, n7979);
  and g14855 (n7980, n1574, n_7516);
  not g14856 (n_7517, n7980);
  and g14857 (n7981, n1576, n_7517);
  not g14858 (n_7518, n7981);
  and g14859 (n7982, n1837, n_7518);
  not g14860 (n_7519, n7982);
  and g14861 (n7983, n1068, n_7519);
  not g14862 (n_7520, n7983);
  and g14863 (n7984, n1072, n_7520);
  not g14864 (n_7521, n7984);
  and g14865 (n7985, n1076, n_7521);
  not g14866 (n_7522, n7985);
  and g14867 (n7986, n1080, n_7522);
  not g14868 (n_7523, n7986);
  and g14869 (n7987, n1084, n_7523);
  not g14870 (n_7524, n7987);
  and g14871 (n7988, n1088, n_7524);
  not g14872 (n_7525, n7988);
  and g14873 (n7989, n1092, n_7525);
  not g14874 (n_7526, n7989);
  and g14875 (n7990, n1096, n_7526);
  not g14876 (n_7527, n7990);
  and g14877 (n7991, n1100, n_7527);
  not g14878 (n_7528, n7991);
  and g14879 (n7992, n1104, n_7528);
  not g14880 (n_7529, n7992);
  and g14881 (n7993, n1108, n_7529);
  not g14882 (n_7530, n7993);
  and g14883 (n7994, n1112, n_7530);
  not g14884 (n_7531, n7994);
  and g14885 (n7995, n1116, n_7531);
  not g14886 (n_7532, n7995);
  and g14887 (n7996, n1120, n_7532);
  not g14888 (n_7533, n7996);
  and g14889 (n7997, n1124, n_7533);
  not g14890 (n_7534, n7997);
  and g14891 (n7998, n1128, n_7534);
  not g14892 (n_7535, n7998);
  and g14893 (n7999, n1132, n_7535);
  not g14894 (n_7536, n7999);
  and g14895 (n8000, n1136, n_7536);
  not g14896 (n_7537, n8000);
  and g14897 (n8001, n1140, n_7537);
  not g14898 (n_7538, n8001);
  and g14899 (n8002, n1144, n_7538);
  not g14900 (n_7539, n8002);
  and g14901 (n8003, n1148, n_7539);
  not g14902 (n_7540, n8003);
  and g14903 (n8004, n1152, n_7540);
  not g14904 (n_7541, n8004);
  and g14905 (n8005, n1156, n_7541);
  not g14906 (n_7542, n8005);
  and g14907 (n8006, n1160, n_7542);
  not g14908 (n_7543, n8006);
  and g14909 (n8007, n1164, n_7543);
  not g14910 (n_7544, n8007);
  and g14911 (n8008, n1168, n_7544);
  not g14912 (n_7545, n8008);
  and g14913 (n8009, n1172, n_7545);
  not g14914 (n_7546, n8009);
  and g14915 (n8010, n1176, n_7546);
  not g14916 (n_7547, n8010);
  and g14917 (n8011, n1180, n_7547);
  not g14918 (n_7548, n8011);
  and g14919 (n8012, n1184, n_7548);
  not g14920 (n_7549, n8012);
  and g14921 (n8013, n1188, n_7549);
  not g14922 (n_7550, n8013);
  and g14923 (n8014, n1192, n_7550);
  not g14924 (n_7551, n8014);
  and g14925 (n8015, n1196, n_7551);
  not g14926 (n_7552, n8015);
  and g14927 (n8016, n1200, n_7552);
  not g14928 (n_7553, n8016);
  and g14929 (n8017, n1204, n_7553);
  not g14930 (n_7554, n8017);
  and g14931 (n8018, n1208, n_7554);
  not g14932 (n_7555, n8018);
  and g14933 (n8019, n1212, n_7555);
  not g14934 (n_7556, n8019);
  and g14935 (n8020, n1216, n_7556);
  not g14936 (n_7557, n8020);
  and g14937 (n8021, n1220, n_7557);
  not g14938 (n_7558, n8021);
  and g14939 (n8022, n1224, n_7558);
  not g14940 (n_7559, n8022);
  and g14941 (n8023, n1228, n_7559);
  not g14942 (n_7560, n8023);
  and g14943 (n8024, n1232, n_7560);
  not g14944 (n_7561, n8024);
  and g14945 (n8025, n1236, n_7561);
  not g14946 (n_7562, n8025);
  and g14947 (n8026, n1240, n_7562);
  not g14948 (n_7563, n8026);
  and g14949 (n8027, n1244, n_7563);
  not g14950 (n_7564, n8027);
  and g14951 (n8028, n1248, n_7564);
  not g14952 (n_7565, n8028);
  and g14953 (n8029, n1252, n_7565);
  not g14954 (n_7566, n8029);
  and g14955 (n8030, n1256, n_7566);
  not g14956 (n_7567, n8030);
  and g14957 (n8031, n1260, n_7567);
  and g14958 (n8032, \req[79] , n_951);
  not g14959 (n_7568, n8031);
  and g14960 (\grant[79] , n_7568, n8032);
  not g14961 (n_7569, n599);
  and g14962 (n8034, n_7569, n1271);
  not g14963 (n_7570, n8034);
  and g14964 (n8035, n1276, n_7570);
  not g14965 (n_7571, n8035);
  and g14966 (n8036, n1280, n_7571);
  not g14967 (n_7572, n8036);
  and g14968 (n8037, n1284, n_7572);
  not g14969 (n_7573, n8037);
  and g14970 (n8038, n1288, n_7573);
  not g14971 (n_7574, n8038);
  and g14972 (n8039, n1292, n_7574);
  not g14973 (n_7575, n8039);
  and g14974 (n8040, n1296, n_7575);
  not g14975 (n_7576, n8040);
  and g14976 (n8041, n1300, n_7576);
  not g14977 (n_7577, n8041);
  and g14978 (n8042, n1304, n_7577);
  not g14979 (n_7578, n8042);
  and g14980 (n8043, n1308, n_7578);
  not g14981 (n_7579, n8043);
  and g14982 (n8044, n1312, n_7579);
  not g14983 (n_7580, n8044);
  and g14984 (n8045, n1316, n_7580);
  not g14985 (n_7581, n8045);
  and g14986 (n8046, n1320, n_7581);
  not g14987 (n_7582, n8046);
  and g14988 (n8047, n1324, n_7582);
  not g14989 (n_7583, n8047);
  and g14990 (n8048, n1328, n_7583);
  not g14991 (n_7584, n8048);
  and g14992 (n8049, n1332, n_7584);
  not g14993 (n_7585, n8049);
  and g14994 (n8050, n1336, n_7585);
  not g14995 (n_7586, n8050);
  and g14996 (n8051, n1340, n_7586);
  not g14997 (n_7587, n8051);
  and g14998 (n8052, n1344, n_7587);
  not g14999 (n_7588, n8052);
  and g15000 (n8053, n1348, n_7588);
  not g15001 (n_7589, n8053);
  and g15002 (n8054, n1352, n_7589);
  not g15003 (n_7590, n8054);
  and g15004 (n8055, n1356, n_7590);
  not g15005 (n_7591, n8055);
  and g15006 (n8056, n1360, n_7591);
  not g15007 (n_7592, n8056);
  and g15008 (n8057, n1364, n_7592);
  not g15009 (n_7593, n8057);
  and g15010 (n8058, n1368, n_7593);
  not g15011 (n_7594, n8058);
  and g15012 (n8059, n1372, n_7594);
  not g15013 (n_7595, n8059);
  and g15014 (n8060, n1376, n_7595);
  not g15015 (n_7596, n8060);
  and g15016 (n8061, n1380, n_7596);
  not g15017 (n_7597, n8061);
  and g15018 (n8062, n1384, n_7597);
  not g15019 (n_7598, n8062);
  and g15020 (n8063, n1388, n_7598);
  not g15021 (n_7599, n8063);
  and g15022 (n8064, n1392, n_7599);
  not g15023 (n_7600, n8064);
  and g15024 (n8065, n1396, n_7600);
  not g15025 (n_7601, n8065);
  and g15026 (n8066, n1663, n_7601);
  not g15027 (n_7602, n8066);
  and g15028 (n8067, n392, n_7602);
  not g15029 (n_7603, n8067);
  and g15030 (n8068, n396, n_7603);
  not g15031 (n_7604, n8068);
  and g15032 (n8069, n400, n_7604);
  not g15033 (n_7605, n8069);
  and g15034 (n8070, n404, n_7605);
  not g15035 (n_7606, n8070);
  and g15036 (n8071, n408, n_7606);
  not g15037 (n_7607, n8071);
  and g15038 (n8072, n412, n_7607);
  not g15039 (n_7608, n8072);
  and g15040 (n8073, n416, n_7608);
  not g15041 (n_7609, n8073);
  and g15042 (n8074, n420, n_7609);
  not g15043 (n_7610, n8074);
  and g15044 (n8075, n424, n_7610);
  not g15045 (n_7611, n8075);
  and g15046 (n8076, n428, n_7611);
  not g15047 (n_7612, n8076);
  and g15048 (n8077, n432, n_7612);
  not g15049 (n_7613, n8077);
  and g15050 (n8078, n436, n_7613);
  not g15051 (n_7614, n8078);
  and g15052 (n8079, n440, n_7614);
  not g15053 (n_7615, n8079);
  and g15054 (n8080, n444, n_7615);
  not g15055 (n_7616, n8080);
  and g15056 (n8081, n448, n_7616);
  not g15057 (n_7617, n8081);
  and g15058 (n8082, n452, n_7617);
  not g15059 (n_7618, n8082);
  and g15060 (n8083, n456, n_7618);
  not g15061 (n_7619, n8083);
  and g15062 (n8084, n460, n_7619);
  not g15063 (n_7620, n8084);
  and g15064 (n8085, n464, n_7620);
  not g15065 (n_7621, n8085);
  and g15066 (n8086, n468, n_7621);
  not g15067 (n_7622, n8086);
  and g15068 (n8087, n472, n_7622);
  not g15069 (n_7623, n8087);
  and g15070 (n8088, n476, n_7623);
  not g15071 (n_7624, n8088);
  and g15072 (n8089, n480, n_7624);
  not g15073 (n_7625, n8089);
  and g15074 (n8090, n484, n_7625);
  not g15075 (n_7626, n8090);
  and g15076 (n8091, n488, n_7626);
  not g15077 (n_7627, n8091);
  and g15078 (n8092, n492, n_7627);
  not g15079 (n_7628, n8092);
  and g15080 (n8093, n496, n_7628);
  not g15081 (n_7629, n8093);
  and g15082 (n8094, n500, n_7629);
  not g15083 (n_7630, n8094);
  and g15084 (n8095, n504, n_7630);
  not g15085 (n_7631, n8095);
  and g15086 (n8096, n508, n_7631);
  not g15087 (n_7632, n8096);
  and g15088 (n8097, n512, n_7632);
  not g15089 (n_7633, n8097);
  and g15090 (n8098, n516, n_7633);
  not g15091 (n_7634, n8098);
  and g15092 (n8099, n520, n_7634);
  not g15093 (n_7635, n8099);
  and g15094 (n8100, n524, n_7635);
  not g15095 (n_7636, n8100);
  and g15096 (n8101, n528, n_7636);
  not g15097 (n_7637, n8101);
  and g15098 (n8102, n532, n_7637);
  not g15099 (n_7638, n8102);
  and g15100 (n8103, n536, n_7638);
  not g15101 (n_7639, n8103);
  and g15102 (n8104, n540, n_7639);
  not g15103 (n_7640, n8104);
  and g15104 (n8105, n544, n_7640);
  not g15105 (n_7641, n8105);
  and g15106 (n8106, n548, n_7641);
  not g15107 (n_7642, n8106);
  and g15108 (n8107, n552, n_7642);
  not g15109 (n_7643, n8107);
  and g15110 (n8108, n556, n_7643);
  not g15111 (n_7644, n8108);
  and g15112 (n8109, n560, n_7644);
  not g15113 (n_7645, n8109);
  and g15114 (n8110, n564, n_7645);
  not g15115 (n_7646, n8110);
  and g15116 (n8111, n568, n_7646);
  not g15117 (n_7647, n8111);
  and g15118 (n8112, n572, n_7647);
  not g15119 (n_7648, n8112);
  and g15120 (n8113, n576, n_7648);
  not g15121 (n_7649, n8113);
  and g15122 (n8114, n580, n_7649);
  not g15123 (n_7650, n8114);
  and g15124 (n8115, n584, n_7650);
  not g15125 (n_7651, n8115);
  and g15126 (n8116, n588, n_7651);
  not g15127 (n_7652, n8116);
  and g15128 (n8117, n592, n_7652);
  and g15129 (n8118, \req[80] , n_374);
  not g15130 (n_7653, n8117);
  and g15131 (\grant[80] , n_7653, n8118);
  not g15132 (n_7654, n938);
  and g15133 (n8120, n603, n_7654);
  not g15134 (n_7655, n8120);
  and g15135 (n8121, n608, n_7655);
  not g15136 (n_7656, n8121);
  and g15137 (n8122, n612, n_7656);
  not g15138 (n_7657, n8122);
  and g15139 (n8123, n616, n_7657);
  not g15140 (n_7658, n8123);
  and g15141 (n8124, n620, n_7658);
  not g15142 (n_7659, n8124);
  and g15143 (n8125, n624, n_7659);
  not g15144 (n_7660, n8125);
  and g15145 (n8126, n628, n_7660);
  not g15146 (n_7661, n8126);
  and g15147 (n8127, n632, n_7661);
  not g15148 (n_7662, n8127);
  and g15149 (n8128, n636, n_7662);
  not g15150 (n_7663, n8128);
  and g15151 (n8129, n640, n_7663);
  not g15152 (n_7664, n8129);
  and g15153 (n8130, n644, n_7664);
  not g15154 (n_7665, n8130);
  and g15155 (n8131, n648, n_7665);
  not g15156 (n_7666, n8131);
  and g15157 (n8132, n652, n_7666);
  not g15158 (n_7667, n8132);
  and g15159 (n8133, n656, n_7667);
  not g15160 (n_7668, n8133);
  and g15161 (n8134, n660, n_7668);
  not g15162 (n_7669, n8134);
  and g15163 (n8135, n664, n_7669);
  not g15164 (n_7670, n8135);
  and g15165 (n8136, n668, n_7670);
  not g15166 (n_7671, n8136);
  and g15167 (n8137, n672, n_7671);
  not g15168 (n_7672, n8137);
  and g15169 (n8138, n676, n_7672);
  not g15170 (n_7673, n8138);
  and g15171 (n8139, n680, n_7673);
  not g15172 (n_7674, n8139);
  and g15173 (n8140, n684, n_7674);
  not g15174 (n_7675, n8140);
  and g15175 (n8141, n688, n_7675);
  not g15176 (n_7676, n8141);
  and g15177 (n8142, n692, n_7676);
  not g15178 (n_7677, n8142);
  and g15179 (n8143, n696, n_7677);
  not g15180 (n_7678, n8143);
  and g15181 (n8144, n700, n_7678);
  not g15182 (n_7679, n8144);
  and g15183 (n8145, n704, n_7679);
  not g15184 (n_7680, n8145);
  and g15185 (n8146, n708, n_7680);
  not g15186 (n_7681, n8146);
  and g15187 (n8147, n712, n_7681);
  not g15188 (n_7682, n8147);
  and g15189 (n8148, n716, n_7682);
  not g15190 (n_7683, n8148);
  and g15191 (n8149, n720, n_7683);
  not g15192 (n_7684, n8149);
  and g15193 (n8150, n1484, n_7684);
  not g15194 (n_7685, n8150);
  and g15195 (n8151, n1486, n_7685);
  not g15196 (n_7686, n8151);
  and g15197 (n8152, n1750, n_7686);
  not g15198 (n_7687, n8152);
  and g15199 (n8153, n731, n_7687);
  not g15200 (n_7688, n8153);
  and g15201 (n8154, n735, n_7688);
  not g15202 (n_7689, n8154);
  and g15203 (n8155, n739, n_7689);
  not g15204 (n_7690, n8155);
  and g15205 (n8156, n743, n_7690);
  not g15206 (n_7691, n8156);
  and g15207 (n8157, n747, n_7691);
  not g15208 (n_7692, n8157);
  and g15209 (n8158, n751, n_7692);
  not g15210 (n_7693, n8158);
  and g15211 (n8159, n755, n_7693);
  not g15212 (n_7694, n8159);
  and g15213 (n8160, n759, n_7694);
  not g15214 (n_7695, n8160);
  and g15215 (n8161, n763, n_7695);
  not g15216 (n_7696, n8161);
  and g15217 (n8162, n767, n_7696);
  not g15218 (n_7697, n8162);
  and g15219 (n8163, n771, n_7697);
  not g15220 (n_7698, n8163);
  and g15221 (n8164, n775, n_7698);
  not g15222 (n_7699, n8164);
  and g15223 (n8165, n779, n_7699);
  not g15224 (n_7700, n8165);
  and g15225 (n8166, n783, n_7700);
  not g15226 (n_7701, n8166);
  and g15227 (n8167, n787, n_7701);
  not g15228 (n_7702, n8167);
  and g15229 (n8168, n791, n_7702);
  not g15230 (n_7703, n8168);
  and g15231 (n8169, n795, n_7703);
  not g15232 (n_7704, n8169);
  and g15233 (n8170, n799, n_7704);
  not g15234 (n_7705, n8170);
  and g15235 (n8171, n803, n_7705);
  not g15236 (n_7706, n8171);
  and g15237 (n8172, n807, n_7706);
  not g15238 (n_7707, n8172);
  and g15239 (n8173, n811, n_7707);
  not g15240 (n_7708, n8173);
  and g15241 (n8174, n815, n_7708);
  not g15242 (n_7709, n8174);
  and g15243 (n8175, n819, n_7709);
  not g15244 (n_7710, n8175);
  and g15245 (n8176, n823, n_7710);
  not g15246 (n_7711, n8176);
  and g15247 (n8177, n827, n_7711);
  not g15248 (n_7712, n8177);
  and g15249 (n8178, n831, n_7712);
  not g15250 (n_7713, n8178);
  and g15251 (n8179, n835, n_7713);
  not g15252 (n_7714, n8179);
  and g15253 (n8180, n839, n_7714);
  not g15254 (n_7715, n8180);
  and g15255 (n8181, n843, n_7715);
  not g15256 (n_7716, n8181);
  and g15257 (n8182, n847, n_7716);
  not g15258 (n_7717, n8182);
  and g15259 (n8183, n851, n_7717);
  not g15260 (n_7718, n8183);
  and g15261 (n8184, n855, n_7718);
  not g15262 (n_7719, n8184);
  and g15263 (n8185, n859, n_7719);
  not g15264 (n_7720, n8185);
  and g15265 (n8186, n863, n_7720);
  not g15266 (n_7721, n8186);
  and g15267 (n8187, n867, n_7721);
  not g15268 (n_7722, n8187);
  and g15269 (n8188, n871, n_7722);
  not g15270 (n_7723, n8188);
  and g15271 (n8189, n875, n_7723);
  not g15272 (n_7724, n8189);
  and g15273 (n8190, n879, n_7724);
  not g15274 (n_7725, n8190);
  and g15275 (n8191, n883, n_7725);
  not g15276 (n_7726, n8191);
  and g15277 (n8192, n887, n_7726);
  not g15278 (n_7727, n8192);
  and g15279 (n8193, n891, n_7727);
  not g15280 (n_7728, n8193);
  and g15281 (n8194, n895, n_7728);
  not g15282 (n_7729, n8194);
  and g15283 (n8195, n899, n_7729);
  not g15284 (n_7730, n8195);
  and g15285 (n8196, n903, n_7730);
  not g15286 (n_7731, n8196);
  and g15287 (n8197, n907, n_7731);
  not g15288 (n_7732, n8197);
  and g15289 (n8198, n911, n_7732);
  not g15290 (n_7733, n8198);
  and g15291 (n8199, n915, n_7733);
  not g15292 (n_7734, n8199);
  and g15293 (n8200, n919, n_7734);
  not g15294 (n_7735, n8200);
  and g15295 (n8201, n923, n_7735);
  not g15296 (n_7736, n8201);
  and g15297 (n8202, n927, n_7736);
  not g15298 (n_7737, n8202);
  and g15299 (n8203, n931, n_7737);
  and g15300 (n8204, \req[81] , n_755);
  not g15301 (n_7738, n8203);
  and g15302 (\grant[81] , n_7738, n8204);
  not g15303 (n_7739, n1275);
  and g15304 (n8206, n942, n_7739);
  not g15305 (n_7740, n8206);
  and g15306 (n8207, n947, n_7740);
  not g15307 (n_7741, n8207);
  and g15308 (n8208, n951, n_7741);
  not g15309 (n_7742, n8208);
  and g15310 (n8209, n955, n_7742);
  not g15311 (n_7743, n8209);
  and g15312 (n8210, n959, n_7743);
  not g15313 (n_7744, n8210);
  and g15314 (n8211, n963, n_7744);
  not g15315 (n_7745, n8211);
  and g15316 (n8212, n967, n_7745);
  not g15317 (n_7746, n8212);
  and g15318 (n8213, n971, n_7746);
  not g15319 (n_7747, n8213);
  and g15320 (n8214, n975, n_7747);
  not g15321 (n_7748, n8214);
  and g15322 (n8215, n979, n_7748);
  not g15323 (n_7749, n8215);
  and g15324 (n8216, n983, n_7749);
  not g15325 (n_7750, n8216);
  and g15326 (n8217, n987, n_7750);
  not g15327 (n_7751, n8217);
  and g15328 (n8218, n991, n_7751);
  not g15329 (n_7752, n8218);
  and g15330 (n8219, n995, n_7752);
  not g15331 (n_7753, n8219);
  and g15332 (n8220, n999, n_7753);
  not g15333 (n_7754, n8220);
  and g15334 (n8221, n1003, n_7754);
  not g15335 (n_7755, n8221);
  and g15336 (n8222, n1007, n_7755);
  not g15337 (n_7756, n8222);
  and g15338 (n8223, n1011, n_7756);
  not g15339 (n_7757, n8223);
  and g15340 (n8224, n1015, n_7757);
  not g15341 (n_7758, n8224);
  and g15342 (n8225, n1019, n_7758);
  not g15343 (n_7759, n8225);
  and g15344 (n8226, n1023, n_7759);
  not g15345 (n_7760, n8226);
  and g15346 (n8227, n1027, n_7760);
  not g15347 (n_7761, n8227);
  and g15348 (n8228, n1031, n_7761);
  not g15349 (n_7762, n8228);
  and g15350 (n8229, n1035, n_7762);
  not g15351 (n_7763, n8229);
  and g15352 (n8230, n1039, n_7763);
  not g15353 (n_7764, n8230);
  and g15354 (n8231, n1043, n_7764);
  not g15355 (n_7765, n8231);
  and g15356 (n8232, n1047, n_7765);
  not g15357 (n_7766, n8232);
  and g15358 (n8233, n1051, n_7766);
  not g15359 (n_7767, n8233);
  and g15360 (n8234, n1055, n_7767);
  not g15361 (n_7768, n8234);
  and g15362 (n8235, n1059, n_7768);
  not g15363 (n_7769, n8235);
  and g15364 (n8236, n1574, n_7769);
  not g15365 (n_7770, n8236);
  and g15366 (n8237, n1576, n_7770);
  not g15367 (n_7771, n8237);
  and g15368 (n8238, n1837, n_7771);
  not g15369 (n_7772, n8238);
  and g15370 (n8239, n1068, n_7772);
  not g15371 (n_7773, n8239);
  and g15372 (n8240, n1072, n_7773);
  not g15373 (n_7774, n8240);
  and g15374 (n8241, n1076, n_7774);
  not g15375 (n_7775, n8241);
  and g15376 (n8242, n1080, n_7775);
  not g15377 (n_7776, n8242);
  and g15378 (n8243, n1084, n_7776);
  not g15379 (n_7777, n8243);
  and g15380 (n8244, n1088, n_7777);
  not g15381 (n_7778, n8244);
  and g15382 (n8245, n1092, n_7778);
  not g15383 (n_7779, n8245);
  and g15384 (n8246, n1096, n_7779);
  not g15385 (n_7780, n8246);
  and g15386 (n8247, n1100, n_7780);
  not g15387 (n_7781, n8247);
  and g15388 (n8248, n1104, n_7781);
  not g15389 (n_7782, n8248);
  and g15390 (n8249, n1108, n_7782);
  not g15391 (n_7783, n8249);
  and g15392 (n8250, n1112, n_7783);
  not g15393 (n_7784, n8250);
  and g15394 (n8251, n1116, n_7784);
  not g15395 (n_7785, n8251);
  and g15396 (n8252, n1120, n_7785);
  not g15397 (n_7786, n8252);
  and g15398 (n8253, n1124, n_7786);
  not g15399 (n_7787, n8253);
  and g15400 (n8254, n1128, n_7787);
  not g15401 (n_7788, n8254);
  and g15402 (n8255, n1132, n_7788);
  not g15403 (n_7789, n8255);
  and g15404 (n8256, n1136, n_7789);
  not g15405 (n_7790, n8256);
  and g15406 (n8257, n1140, n_7790);
  not g15407 (n_7791, n8257);
  and g15408 (n8258, n1144, n_7791);
  not g15409 (n_7792, n8258);
  and g15410 (n8259, n1148, n_7792);
  not g15411 (n_7793, n8259);
  and g15412 (n8260, n1152, n_7793);
  not g15413 (n_7794, n8260);
  and g15414 (n8261, n1156, n_7794);
  not g15415 (n_7795, n8261);
  and g15416 (n8262, n1160, n_7795);
  not g15417 (n_7796, n8262);
  and g15418 (n8263, n1164, n_7796);
  not g15419 (n_7797, n8263);
  and g15420 (n8264, n1168, n_7797);
  not g15421 (n_7798, n8264);
  and g15422 (n8265, n1172, n_7798);
  not g15423 (n_7799, n8265);
  and g15424 (n8266, n1176, n_7799);
  not g15425 (n_7800, n8266);
  and g15426 (n8267, n1180, n_7800);
  not g15427 (n_7801, n8267);
  and g15428 (n8268, n1184, n_7801);
  not g15429 (n_7802, n8268);
  and g15430 (n8269, n1188, n_7802);
  not g15431 (n_7803, n8269);
  and g15432 (n8270, n1192, n_7803);
  not g15433 (n_7804, n8270);
  and g15434 (n8271, n1196, n_7804);
  not g15435 (n_7805, n8271);
  and g15436 (n8272, n1200, n_7805);
  not g15437 (n_7806, n8272);
  and g15438 (n8273, n1204, n_7806);
  not g15439 (n_7807, n8273);
  and g15440 (n8274, n1208, n_7807);
  not g15441 (n_7808, n8274);
  and g15442 (n8275, n1212, n_7808);
  not g15443 (n_7809, n8275);
  and g15444 (n8276, n1216, n_7809);
  not g15445 (n_7810, n8276);
  and g15446 (n8277, n1220, n_7810);
  not g15447 (n_7811, n8277);
  and g15448 (n8278, n1224, n_7811);
  not g15449 (n_7812, n8278);
  and g15450 (n8279, n1228, n_7812);
  not g15451 (n_7813, n8279);
  and g15452 (n8280, n1232, n_7813);
  not g15453 (n_7814, n8280);
  and g15454 (n8281, n1236, n_7814);
  not g15455 (n_7815, n8281);
  and g15456 (n8282, n1240, n_7815);
  not g15457 (n_7816, n8282);
  and g15458 (n8283, n1244, n_7816);
  not g15459 (n_7817, n8283);
  and g15460 (n8284, n1248, n_7817);
  not g15461 (n_7818, n8284);
  and g15462 (n8285, n1252, n_7818);
  not g15463 (n_7819, n8285);
  and g15464 (n8286, n1256, n_7819);
  not g15465 (n_7820, n8286);
  and g15466 (n8287, n1260, n_7820);
  not g15467 (n_7821, n8287);
  and g15468 (n8288, n1264, n_7821);
  not g15469 (n_7822, n8288);
  and g15470 (n8289, n1268, n_7822);
  and g15471 (n8290, \req[82] , n_955);
  not g15472 (n_7823, n8289);
  and g15473 (\grant[82] , n_7823, n8290);
  not g15474 (n_7824, n607);
  and g15475 (n8292, n_7824, n1279);
  not g15476 (n_7825, n8292);
  and g15477 (n8293, n1284, n_7825);
  not g15478 (n_7826, n8293);
  and g15479 (n8294, n1288, n_7826);
  not g15480 (n_7827, n8294);
  and g15481 (n8295, n1292, n_7827);
  not g15482 (n_7828, n8295);
  and g15483 (n8296, n1296, n_7828);
  not g15484 (n_7829, n8296);
  and g15485 (n8297, n1300, n_7829);
  not g15486 (n_7830, n8297);
  and g15487 (n8298, n1304, n_7830);
  not g15488 (n_7831, n8298);
  and g15489 (n8299, n1308, n_7831);
  not g15490 (n_7832, n8299);
  and g15491 (n8300, n1312, n_7832);
  not g15492 (n_7833, n8300);
  and g15493 (n8301, n1316, n_7833);
  not g15494 (n_7834, n8301);
  and g15495 (n8302, n1320, n_7834);
  not g15496 (n_7835, n8302);
  and g15497 (n8303, n1324, n_7835);
  not g15498 (n_7836, n8303);
  and g15499 (n8304, n1328, n_7836);
  not g15500 (n_7837, n8304);
  and g15501 (n8305, n1332, n_7837);
  not g15502 (n_7838, n8305);
  and g15503 (n8306, n1336, n_7838);
  not g15504 (n_7839, n8306);
  and g15505 (n8307, n1340, n_7839);
  not g15506 (n_7840, n8307);
  and g15507 (n8308, n1344, n_7840);
  not g15508 (n_7841, n8308);
  and g15509 (n8309, n1348, n_7841);
  not g15510 (n_7842, n8309);
  and g15511 (n8310, n1352, n_7842);
  not g15512 (n_7843, n8310);
  and g15513 (n8311, n1356, n_7843);
  not g15514 (n_7844, n8311);
  and g15515 (n8312, n1360, n_7844);
  not g15516 (n_7845, n8312);
  and g15517 (n8313, n1364, n_7845);
  not g15518 (n_7846, n8313);
  and g15519 (n8314, n1368, n_7846);
  not g15520 (n_7847, n8314);
  and g15521 (n8315, n1372, n_7847);
  not g15522 (n_7848, n8315);
  and g15523 (n8316, n1376, n_7848);
  not g15524 (n_7849, n8316);
  and g15525 (n8317, n1380, n_7849);
  not g15526 (n_7850, n8317);
  and g15527 (n8318, n1384, n_7850);
  not g15528 (n_7851, n8318);
  and g15529 (n8319, n1388, n_7851);
  not g15530 (n_7852, n8319);
  and g15531 (n8320, n1392, n_7852);
  not g15532 (n_7853, n8320);
  and g15533 (n8321, n1396, n_7853);
  not g15534 (n_7854, n8321);
  and g15535 (n8322, n1663, n_7854);
  not g15536 (n_7855, n8322);
  and g15537 (n8323, n392, n_7855);
  not g15538 (n_7856, n8323);
  and g15539 (n8324, n396, n_7856);
  not g15540 (n_7857, n8324);
  and g15541 (n8325, n400, n_7857);
  not g15542 (n_7858, n8325);
  and g15543 (n8326, n404, n_7858);
  not g15544 (n_7859, n8326);
  and g15545 (n8327, n408, n_7859);
  not g15546 (n_7860, n8327);
  and g15547 (n8328, n412, n_7860);
  not g15548 (n_7861, n8328);
  and g15549 (n8329, n416, n_7861);
  not g15550 (n_7862, n8329);
  and g15551 (n8330, n420, n_7862);
  not g15552 (n_7863, n8330);
  and g15553 (n8331, n424, n_7863);
  not g15554 (n_7864, n8331);
  and g15555 (n8332, n428, n_7864);
  not g15556 (n_7865, n8332);
  and g15557 (n8333, n432, n_7865);
  not g15558 (n_7866, n8333);
  and g15559 (n8334, n436, n_7866);
  not g15560 (n_7867, n8334);
  and g15561 (n8335, n440, n_7867);
  not g15562 (n_7868, n8335);
  and g15563 (n8336, n444, n_7868);
  not g15564 (n_7869, n8336);
  and g15565 (n8337, n448, n_7869);
  not g15566 (n_7870, n8337);
  and g15567 (n8338, n452, n_7870);
  not g15568 (n_7871, n8338);
  and g15569 (n8339, n456, n_7871);
  not g15570 (n_7872, n8339);
  and g15571 (n8340, n460, n_7872);
  not g15572 (n_7873, n8340);
  and g15573 (n8341, n464, n_7873);
  not g15574 (n_7874, n8341);
  and g15575 (n8342, n468, n_7874);
  not g15576 (n_7875, n8342);
  and g15577 (n8343, n472, n_7875);
  not g15578 (n_7876, n8343);
  and g15579 (n8344, n476, n_7876);
  not g15580 (n_7877, n8344);
  and g15581 (n8345, n480, n_7877);
  not g15582 (n_7878, n8345);
  and g15583 (n8346, n484, n_7878);
  not g15584 (n_7879, n8346);
  and g15585 (n8347, n488, n_7879);
  not g15586 (n_7880, n8347);
  and g15587 (n8348, n492, n_7880);
  not g15588 (n_7881, n8348);
  and g15589 (n8349, n496, n_7881);
  not g15590 (n_7882, n8349);
  and g15591 (n8350, n500, n_7882);
  not g15592 (n_7883, n8350);
  and g15593 (n8351, n504, n_7883);
  not g15594 (n_7884, n8351);
  and g15595 (n8352, n508, n_7884);
  not g15596 (n_7885, n8352);
  and g15597 (n8353, n512, n_7885);
  not g15598 (n_7886, n8353);
  and g15599 (n8354, n516, n_7886);
  not g15600 (n_7887, n8354);
  and g15601 (n8355, n520, n_7887);
  not g15602 (n_7888, n8355);
  and g15603 (n8356, n524, n_7888);
  not g15604 (n_7889, n8356);
  and g15605 (n8357, n528, n_7889);
  not g15606 (n_7890, n8357);
  and g15607 (n8358, n532, n_7890);
  not g15608 (n_7891, n8358);
  and g15609 (n8359, n536, n_7891);
  not g15610 (n_7892, n8359);
  and g15611 (n8360, n540, n_7892);
  not g15612 (n_7893, n8360);
  and g15613 (n8361, n544, n_7893);
  not g15614 (n_7894, n8361);
  and g15615 (n8362, n548, n_7894);
  not g15616 (n_7895, n8362);
  and g15617 (n8363, n552, n_7895);
  not g15618 (n_7896, n8363);
  and g15619 (n8364, n556, n_7896);
  not g15620 (n_7897, n8364);
  and g15621 (n8365, n560, n_7897);
  not g15622 (n_7898, n8365);
  and g15623 (n8366, n564, n_7898);
  not g15624 (n_7899, n8366);
  and g15625 (n8367, n568, n_7899);
  not g15626 (n_7900, n8367);
  and g15627 (n8368, n572, n_7900);
  not g15628 (n_7901, n8368);
  and g15629 (n8369, n576, n_7901);
  not g15630 (n_7902, n8369);
  and g15631 (n8370, n580, n_7902);
  not g15632 (n_7903, n8370);
  and g15633 (n8371, n584, n_7903);
  not g15634 (n_7904, n8371);
  and g15635 (n8372, n588, n_7904);
  not g15636 (n_7905, n8372);
  and g15637 (n8373, n592, n_7905);
  not g15638 (n_7906, n8373);
  and g15639 (n8374, n596, n_7906);
  not g15640 (n_7907, n8374);
  and g15641 (n8375, n600, n_7907);
  and g15642 (n8376, \req[83] , n_388);
  not g15643 (n_7908, n8375);
  and g15644 (\grant[83] , n_7908, n8376);
  not g15645 (n_7909, n946);
  and g15646 (n8378, n611, n_7909);
  not g15647 (n_7910, n8378);
  and g15648 (n8379, n616, n_7910);
  not g15649 (n_7911, n8379);
  and g15650 (n8380, n620, n_7911);
  not g15651 (n_7912, n8380);
  and g15652 (n8381, n624, n_7912);
  not g15653 (n_7913, n8381);
  and g15654 (n8382, n628, n_7913);
  not g15655 (n_7914, n8382);
  and g15656 (n8383, n632, n_7914);
  not g15657 (n_7915, n8383);
  and g15658 (n8384, n636, n_7915);
  not g15659 (n_7916, n8384);
  and g15660 (n8385, n640, n_7916);
  not g15661 (n_7917, n8385);
  and g15662 (n8386, n644, n_7917);
  not g15663 (n_7918, n8386);
  and g15664 (n8387, n648, n_7918);
  not g15665 (n_7919, n8387);
  and g15666 (n8388, n652, n_7919);
  not g15667 (n_7920, n8388);
  and g15668 (n8389, n656, n_7920);
  not g15669 (n_7921, n8389);
  and g15670 (n8390, n660, n_7921);
  not g15671 (n_7922, n8390);
  and g15672 (n8391, n664, n_7922);
  not g15673 (n_7923, n8391);
  and g15674 (n8392, n668, n_7923);
  not g15675 (n_7924, n8392);
  and g15676 (n8393, n672, n_7924);
  not g15677 (n_7925, n8393);
  and g15678 (n8394, n676, n_7925);
  not g15679 (n_7926, n8394);
  and g15680 (n8395, n680, n_7926);
  not g15681 (n_7927, n8395);
  and g15682 (n8396, n684, n_7927);
  not g15683 (n_7928, n8396);
  and g15684 (n8397, n688, n_7928);
  not g15685 (n_7929, n8397);
  and g15686 (n8398, n692, n_7929);
  not g15687 (n_7930, n8398);
  and g15688 (n8399, n696, n_7930);
  not g15689 (n_7931, n8399);
  and g15690 (n8400, n700, n_7931);
  not g15691 (n_7932, n8400);
  and g15692 (n8401, n704, n_7932);
  not g15693 (n_7933, n8401);
  and g15694 (n8402, n708, n_7933);
  not g15695 (n_7934, n8402);
  and g15696 (n8403, n712, n_7934);
  not g15697 (n_7935, n8403);
  and g15698 (n8404, n716, n_7935);
  not g15699 (n_7936, n8404);
  and g15700 (n8405, n720, n_7936);
  not g15701 (n_7937, n8405);
  and g15702 (n8406, n1484, n_7937);
  not g15703 (n_7938, n8406);
  and g15704 (n8407, n1486, n_7938);
  not g15705 (n_7939, n8407);
  and g15706 (n8408, n1750, n_7939);
  not g15707 (n_7940, n8408);
  and g15708 (n8409, n731, n_7940);
  not g15709 (n_7941, n8409);
  and g15710 (n8410, n735, n_7941);
  not g15711 (n_7942, n8410);
  and g15712 (n8411, n739, n_7942);
  not g15713 (n_7943, n8411);
  and g15714 (n8412, n743, n_7943);
  not g15715 (n_7944, n8412);
  and g15716 (n8413, n747, n_7944);
  not g15717 (n_7945, n8413);
  and g15718 (n8414, n751, n_7945);
  not g15719 (n_7946, n8414);
  and g15720 (n8415, n755, n_7946);
  not g15721 (n_7947, n8415);
  and g15722 (n8416, n759, n_7947);
  not g15723 (n_7948, n8416);
  and g15724 (n8417, n763, n_7948);
  not g15725 (n_7949, n8417);
  and g15726 (n8418, n767, n_7949);
  not g15727 (n_7950, n8418);
  and g15728 (n8419, n771, n_7950);
  not g15729 (n_7951, n8419);
  and g15730 (n8420, n775, n_7951);
  not g15731 (n_7952, n8420);
  and g15732 (n8421, n779, n_7952);
  not g15733 (n_7953, n8421);
  and g15734 (n8422, n783, n_7953);
  not g15735 (n_7954, n8422);
  and g15736 (n8423, n787, n_7954);
  not g15737 (n_7955, n8423);
  and g15738 (n8424, n791, n_7955);
  not g15739 (n_7956, n8424);
  and g15740 (n8425, n795, n_7956);
  not g15741 (n_7957, n8425);
  and g15742 (n8426, n799, n_7957);
  not g15743 (n_7958, n8426);
  and g15744 (n8427, n803, n_7958);
  not g15745 (n_7959, n8427);
  and g15746 (n8428, n807, n_7959);
  not g15747 (n_7960, n8428);
  and g15748 (n8429, n811, n_7960);
  not g15749 (n_7961, n8429);
  and g15750 (n8430, n815, n_7961);
  not g15751 (n_7962, n8430);
  and g15752 (n8431, n819, n_7962);
  not g15753 (n_7963, n8431);
  and g15754 (n8432, n823, n_7963);
  not g15755 (n_7964, n8432);
  and g15756 (n8433, n827, n_7964);
  not g15757 (n_7965, n8433);
  and g15758 (n8434, n831, n_7965);
  not g15759 (n_7966, n8434);
  and g15760 (n8435, n835, n_7966);
  not g15761 (n_7967, n8435);
  and g15762 (n8436, n839, n_7967);
  not g15763 (n_7968, n8436);
  and g15764 (n8437, n843, n_7968);
  not g15765 (n_7969, n8437);
  and g15766 (n8438, n847, n_7969);
  not g15767 (n_7970, n8438);
  and g15768 (n8439, n851, n_7970);
  not g15769 (n_7971, n8439);
  and g15770 (n8440, n855, n_7971);
  not g15771 (n_7972, n8440);
  and g15772 (n8441, n859, n_7972);
  not g15773 (n_7973, n8441);
  and g15774 (n8442, n863, n_7973);
  not g15775 (n_7974, n8442);
  and g15776 (n8443, n867, n_7974);
  not g15777 (n_7975, n8443);
  and g15778 (n8444, n871, n_7975);
  not g15779 (n_7976, n8444);
  and g15780 (n8445, n875, n_7976);
  not g15781 (n_7977, n8445);
  and g15782 (n8446, n879, n_7977);
  not g15783 (n_7978, n8446);
  and g15784 (n8447, n883, n_7978);
  not g15785 (n_7979, n8447);
  and g15786 (n8448, n887, n_7979);
  not g15787 (n_7980, n8448);
  and g15788 (n8449, n891, n_7980);
  not g15789 (n_7981, n8449);
  and g15790 (n8450, n895, n_7981);
  not g15791 (n_7982, n8450);
  and g15792 (n8451, n899, n_7982);
  not g15793 (n_7983, n8451);
  and g15794 (n8452, n903, n_7983);
  not g15795 (n_7984, n8452);
  and g15796 (n8453, n907, n_7984);
  not g15797 (n_7985, n8453);
  and g15798 (n8454, n911, n_7985);
  not g15799 (n_7986, n8454);
  and g15800 (n8455, n915, n_7986);
  not g15801 (n_7987, n8455);
  and g15802 (n8456, n919, n_7987);
  not g15803 (n_7988, n8456);
  and g15804 (n8457, n923, n_7988);
  not g15805 (n_7989, n8457);
  and g15806 (n8458, n927, n_7989);
  not g15807 (n_7990, n8458);
  and g15808 (n8459, n931, n_7990);
  not g15809 (n_7991, n8459);
  and g15810 (n8460, n935, n_7991);
  not g15811 (n_7992, n8460);
  and g15812 (n8461, n939, n_7992);
  and g15813 (n8462, \req[84] , n_761);
  not g15814 (n_7993, n8461);
  and g15815 (\grant[84] , n_7993, n8462);
  not g15816 (n_7994, n1283);
  and g15817 (n8464, n950, n_7994);
  not g15818 (n_7995, n8464);
  and g15819 (n8465, n955, n_7995);
  not g15820 (n_7996, n8465);
  and g15821 (n8466, n959, n_7996);
  not g15822 (n_7997, n8466);
  and g15823 (n8467, n963, n_7997);
  not g15824 (n_7998, n8467);
  and g15825 (n8468, n967, n_7998);
  not g15826 (n_7999, n8468);
  and g15827 (n8469, n971, n_7999);
  not g15828 (n_8000, n8469);
  and g15829 (n8470, n975, n_8000);
  not g15830 (n_8001, n8470);
  and g15831 (n8471, n979, n_8001);
  not g15832 (n_8002, n8471);
  and g15833 (n8472, n983, n_8002);
  not g15834 (n_8003, n8472);
  and g15835 (n8473, n987, n_8003);
  not g15836 (n_8004, n8473);
  and g15837 (n8474, n991, n_8004);
  not g15838 (n_8005, n8474);
  and g15839 (n8475, n995, n_8005);
  not g15840 (n_8006, n8475);
  and g15841 (n8476, n999, n_8006);
  not g15842 (n_8007, n8476);
  and g15843 (n8477, n1003, n_8007);
  not g15844 (n_8008, n8477);
  and g15845 (n8478, n1007, n_8008);
  not g15846 (n_8009, n8478);
  and g15847 (n8479, n1011, n_8009);
  not g15848 (n_8010, n8479);
  and g15849 (n8480, n1015, n_8010);
  not g15850 (n_8011, n8480);
  and g15851 (n8481, n1019, n_8011);
  not g15852 (n_8012, n8481);
  and g15853 (n8482, n1023, n_8012);
  not g15854 (n_8013, n8482);
  and g15855 (n8483, n1027, n_8013);
  not g15856 (n_8014, n8483);
  and g15857 (n8484, n1031, n_8014);
  not g15858 (n_8015, n8484);
  and g15859 (n8485, n1035, n_8015);
  not g15860 (n_8016, n8485);
  and g15861 (n8486, n1039, n_8016);
  not g15862 (n_8017, n8486);
  and g15863 (n8487, n1043, n_8017);
  not g15864 (n_8018, n8487);
  and g15865 (n8488, n1047, n_8018);
  not g15866 (n_8019, n8488);
  and g15867 (n8489, n1051, n_8019);
  not g15868 (n_8020, n8489);
  and g15869 (n8490, n1055, n_8020);
  not g15870 (n_8021, n8490);
  and g15871 (n8491, n1059, n_8021);
  not g15872 (n_8022, n8491);
  and g15873 (n8492, n1574, n_8022);
  not g15874 (n_8023, n8492);
  and g15875 (n8493, n1576, n_8023);
  not g15876 (n_8024, n8493);
  and g15877 (n8494, n1837, n_8024);
  not g15878 (n_8025, n8494);
  and g15879 (n8495, n1068, n_8025);
  not g15880 (n_8026, n8495);
  and g15881 (n8496, n1072, n_8026);
  not g15882 (n_8027, n8496);
  and g15883 (n8497, n1076, n_8027);
  not g15884 (n_8028, n8497);
  and g15885 (n8498, n1080, n_8028);
  not g15886 (n_8029, n8498);
  and g15887 (n8499, n1084, n_8029);
  not g15888 (n_8030, n8499);
  and g15889 (n8500, n1088, n_8030);
  not g15890 (n_8031, n8500);
  and g15891 (n8501, n1092, n_8031);
  not g15892 (n_8032, n8501);
  and g15893 (n8502, n1096, n_8032);
  not g15894 (n_8033, n8502);
  and g15895 (n8503, n1100, n_8033);
  not g15896 (n_8034, n8503);
  and g15897 (n8504, n1104, n_8034);
  not g15898 (n_8035, n8504);
  and g15899 (n8505, n1108, n_8035);
  not g15900 (n_8036, n8505);
  and g15901 (n8506, n1112, n_8036);
  not g15902 (n_8037, n8506);
  and g15903 (n8507, n1116, n_8037);
  not g15904 (n_8038, n8507);
  and g15905 (n8508, n1120, n_8038);
  not g15906 (n_8039, n8508);
  and g15907 (n8509, n1124, n_8039);
  not g15908 (n_8040, n8509);
  and g15909 (n8510, n1128, n_8040);
  not g15910 (n_8041, n8510);
  and g15911 (n8511, n1132, n_8041);
  not g15912 (n_8042, n8511);
  and g15913 (n8512, n1136, n_8042);
  not g15914 (n_8043, n8512);
  and g15915 (n8513, n1140, n_8043);
  not g15916 (n_8044, n8513);
  and g15917 (n8514, n1144, n_8044);
  not g15918 (n_8045, n8514);
  and g15919 (n8515, n1148, n_8045);
  not g15920 (n_8046, n8515);
  and g15921 (n8516, n1152, n_8046);
  not g15922 (n_8047, n8516);
  and g15923 (n8517, n1156, n_8047);
  not g15924 (n_8048, n8517);
  and g15925 (n8518, n1160, n_8048);
  not g15926 (n_8049, n8518);
  and g15927 (n8519, n1164, n_8049);
  not g15928 (n_8050, n8519);
  and g15929 (n8520, n1168, n_8050);
  not g15930 (n_8051, n8520);
  and g15931 (n8521, n1172, n_8051);
  not g15932 (n_8052, n8521);
  and g15933 (n8522, n1176, n_8052);
  not g15934 (n_8053, n8522);
  and g15935 (n8523, n1180, n_8053);
  not g15936 (n_8054, n8523);
  and g15937 (n8524, n1184, n_8054);
  not g15938 (n_8055, n8524);
  and g15939 (n8525, n1188, n_8055);
  not g15940 (n_8056, n8525);
  and g15941 (n8526, n1192, n_8056);
  not g15942 (n_8057, n8526);
  and g15943 (n8527, n1196, n_8057);
  not g15944 (n_8058, n8527);
  and g15945 (n8528, n1200, n_8058);
  not g15946 (n_8059, n8528);
  and g15947 (n8529, n1204, n_8059);
  not g15948 (n_8060, n8529);
  and g15949 (n8530, n1208, n_8060);
  not g15950 (n_8061, n8530);
  and g15951 (n8531, n1212, n_8061);
  not g15952 (n_8062, n8531);
  and g15953 (n8532, n1216, n_8062);
  not g15954 (n_8063, n8532);
  and g15955 (n8533, n1220, n_8063);
  not g15956 (n_8064, n8533);
  and g15957 (n8534, n1224, n_8064);
  not g15958 (n_8065, n8534);
  and g15959 (n8535, n1228, n_8065);
  not g15960 (n_8066, n8535);
  and g15961 (n8536, n1232, n_8066);
  not g15962 (n_8067, n8536);
  and g15963 (n8537, n1236, n_8067);
  not g15964 (n_8068, n8537);
  and g15965 (n8538, n1240, n_8068);
  not g15966 (n_8069, n8538);
  and g15967 (n8539, n1244, n_8069);
  not g15968 (n_8070, n8539);
  and g15969 (n8540, n1248, n_8070);
  not g15970 (n_8071, n8540);
  and g15971 (n8541, n1252, n_8071);
  not g15972 (n_8072, n8541);
  and g15973 (n8542, n1256, n_8072);
  not g15974 (n_8073, n8542);
  and g15975 (n8543, n1260, n_8073);
  not g15976 (n_8074, n8543);
  and g15977 (n8544, n1264, n_8074);
  not g15978 (n_8075, n8544);
  and g15979 (n8545, n1268, n_8075);
  not g15980 (n_8076, n8545);
  and g15981 (n8546, n1272, n_8076);
  not g15982 (n_8077, n8546);
  and g15983 (n8547, n1276, n_8077);
  and g15984 (n8548, \req[85] , n_959);
  not g15985 (n_8078, n8547);
  and g15986 (\grant[85] , n_8078, n8548);
  not g15987 (n_8079, n615);
  and g15988 (n8550, n_8079, n1287);
  not g15989 (n_8080, n8550);
  and g15990 (n8551, n1292, n_8080);
  not g15991 (n_8081, n8551);
  and g15992 (n8552, n1296, n_8081);
  not g15993 (n_8082, n8552);
  and g15994 (n8553, n1300, n_8082);
  not g15995 (n_8083, n8553);
  and g15996 (n8554, n1304, n_8083);
  not g15997 (n_8084, n8554);
  and g15998 (n8555, n1308, n_8084);
  not g15999 (n_8085, n8555);
  and g16000 (n8556, n1312, n_8085);
  not g16001 (n_8086, n8556);
  and g16002 (n8557, n1316, n_8086);
  not g16003 (n_8087, n8557);
  and g16004 (n8558, n1320, n_8087);
  not g16005 (n_8088, n8558);
  and g16006 (n8559, n1324, n_8088);
  not g16007 (n_8089, n8559);
  and g16008 (n8560, n1328, n_8089);
  not g16009 (n_8090, n8560);
  and g16010 (n8561, n1332, n_8090);
  not g16011 (n_8091, n8561);
  and g16012 (n8562, n1336, n_8091);
  not g16013 (n_8092, n8562);
  and g16014 (n8563, n1340, n_8092);
  not g16015 (n_8093, n8563);
  and g16016 (n8564, n1344, n_8093);
  not g16017 (n_8094, n8564);
  and g16018 (n8565, n1348, n_8094);
  not g16019 (n_8095, n8565);
  and g16020 (n8566, n1352, n_8095);
  not g16021 (n_8096, n8566);
  and g16022 (n8567, n1356, n_8096);
  not g16023 (n_8097, n8567);
  and g16024 (n8568, n1360, n_8097);
  not g16025 (n_8098, n8568);
  and g16026 (n8569, n1364, n_8098);
  not g16027 (n_8099, n8569);
  and g16028 (n8570, n1368, n_8099);
  not g16029 (n_8100, n8570);
  and g16030 (n8571, n1372, n_8100);
  not g16031 (n_8101, n8571);
  and g16032 (n8572, n1376, n_8101);
  not g16033 (n_8102, n8572);
  and g16034 (n8573, n1380, n_8102);
  not g16035 (n_8103, n8573);
  and g16036 (n8574, n1384, n_8103);
  not g16037 (n_8104, n8574);
  and g16038 (n8575, n1388, n_8104);
  not g16039 (n_8105, n8575);
  and g16040 (n8576, n1392, n_8105);
  not g16041 (n_8106, n8576);
  and g16042 (n8577, n1396, n_8106);
  not g16043 (n_8107, n8577);
  and g16044 (n8578, n1663, n_8107);
  not g16045 (n_8108, n8578);
  and g16046 (n8579, n392, n_8108);
  not g16047 (n_8109, n8579);
  and g16048 (n8580, n396, n_8109);
  not g16049 (n_8110, n8580);
  and g16050 (n8581, n400, n_8110);
  not g16051 (n_8111, n8581);
  and g16052 (n8582, n404, n_8111);
  not g16053 (n_8112, n8582);
  and g16054 (n8583, n408, n_8112);
  not g16055 (n_8113, n8583);
  and g16056 (n8584, n412, n_8113);
  not g16057 (n_8114, n8584);
  and g16058 (n8585, n416, n_8114);
  not g16059 (n_8115, n8585);
  and g16060 (n8586, n420, n_8115);
  not g16061 (n_8116, n8586);
  and g16062 (n8587, n424, n_8116);
  not g16063 (n_8117, n8587);
  and g16064 (n8588, n428, n_8117);
  not g16065 (n_8118, n8588);
  and g16066 (n8589, n432, n_8118);
  not g16067 (n_8119, n8589);
  and g16068 (n8590, n436, n_8119);
  not g16069 (n_8120, n8590);
  and g16070 (n8591, n440, n_8120);
  not g16071 (n_8121, n8591);
  and g16072 (n8592, n444, n_8121);
  not g16073 (n_8122, n8592);
  and g16074 (n8593, n448, n_8122);
  not g16075 (n_8123, n8593);
  and g16076 (n8594, n452, n_8123);
  not g16077 (n_8124, n8594);
  and g16078 (n8595, n456, n_8124);
  not g16079 (n_8125, n8595);
  and g16080 (n8596, n460, n_8125);
  not g16081 (n_8126, n8596);
  and g16082 (n8597, n464, n_8126);
  not g16083 (n_8127, n8597);
  and g16084 (n8598, n468, n_8127);
  not g16085 (n_8128, n8598);
  and g16086 (n8599, n472, n_8128);
  not g16087 (n_8129, n8599);
  and g16088 (n8600, n476, n_8129);
  not g16089 (n_8130, n8600);
  and g16090 (n8601, n480, n_8130);
  not g16091 (n_8131, n8601);
  and g16092 (n8602, n484, n_8131);
  not g16093 (n_8132, n8602);
  and g16094 (n8603, n488, n_8132);
  not g16095 (n_8133, n8603);
  and g16096 (n8604, n492, n_8133);
  not g16097 (n_8134, n8604);
  and g16098 (n8605, n496, n_8134);
  not g16099 (n_8135, n8605);
  and g16100 (n8606, n500, n_8135);
  not g16101 (n_8136, n8606);
  and g16102 (n8607, n504, n_8136);
  not g16103 (n_8137, n8607);
  and g16104 (n8608, n508, n_8137);
  not g16105 (n_8138, n8608);
  and g16106 (n8609, n512, n_8138);
  not g16107 (n_8139, n8609);
  and g16108 (n8610, n516, n_8139);
  not g16109 (n_8140, n8610);
  and g16110 (n8611, n520, n_8140);
  not g16111 (n_8141, n8611);
  and g16112 (n8612, n524, n_8141);
  not g16113 (n_8142, n8612);
  and g16114 (n8613, n528, n_8142);
  not g16115 (n_8143, n8613);
  and g16116 (n8614, n532, n_8143);
  not g16117 (n_8144, n8614);
  and g16118 (n8615, n536, n_8144);
  not g16119 (n_8145, n8615);
  and g16120 (n8616, n540, n_8145);
  not g16121 (n_8146, n8616);
  and g16122 (n8617, n544, n_8146);
  not g16123 (n_8147, n8617);
  and g16124 (n8618, n548, n_8147);
  not g16125 (n_8148, n8618);
  and g16126 (n8619, n552, n_8148);
  not g16127 (n_8149, n8619);
  and g16128 (n8620, n556, n_8149);
  not g16129 (n_8150, n8620);
  and g16130 (n8621, n560, n_8150);
  not g16131 (n_8151, n8621);
  and g16132 (n8622, n564, n_8151);
  not g16133 (n_8152, n8622);
  and g16134 (n8623, n568, n_8152);
  not g16135 (n_8153, n8623);
  and g16136 (n8624, n572, n_8153);
  not g16137 (n_8154, n8624);
  and g16138 (n8625, n576, n_8154);
  not g16139 (n_8155, n8625);
  and g16140 (n8626, n580, n_8155);
  not g16141 (n_8156, n8626);
  and g16142 (n8627, n584, n_8156);
  not g16143 (n_8157, n8627);
  and g16144 (n8628, n588, n_8157);
  not g16145 (n_8158, n8628);
  and g16146 (n8629, n592, n_8158);
  not g16147 (n_8159, n8629);
  and g16148 (n8630, n596, n_8159);
  not g16149 (n_8160, n8630);
  and g16150 (n8631, n600, n_8160);
  not g16151 (n_8161, n8631);
  and g16152 (n8632, n604, n_8161);
  not g16153 (n_8162, n8632);
  and g16154 (n8633, n608, n_8162);
  and g16155 (n8634, \req[86] , n_402);
  not g16156 (n_8163, n8633);
  and g16157 (\grant[86] , n_8163, n8634);
  not g16158 (n_8164, n954);
  and g16159 (n8636, n619, n_8164);
  not g16160 (n_8165, n8636);
  and g16161 (n8637, n624, n_8165);
  not g16162 (n_8166, n8637);
  and g16163 (n8638, n628, n_8166);
  not g16164 (n_8167, n8638);
  and g16165 (n8639, n632, n_8167);
  not g16166 (n_8168, n8639);
  and g16167 (n8640, n636, n_8168);
  not g16168 (n_8169, n8640);
  and g16169 (n8641, n640, n_8169);
  not g16170 (n_8170, n8641);
  and g16171 (n8642, n644, n_8170);
  not g16172 (n_8171, n8642);
  and g16173 (n8643, n648, n_8171);
  not g16174 (n_8172, n8643);
  and g16175 (n8644, n652, n_8172);
  not g16176 (n_8173, n8644);
  and g16177 (n8645, n656, n_8173);
  not g16178 (n_8174, n8645);
  and g16179 (n8646, n660, n_8174);
  not g16180 (n_8175, n8646);
  and g16181 (n8647, n664, n_8175);
  not g16182 (n_8176, n8647);
  and g16183 (n8648, n668, n_8176);
  not g16184 (n_8177, n8648);
  and g16185 (n8649, n672, n_8177);
  not g16186 (n_8178, n8649);
  and g16187 (n8650, n676, n_8178);
  not g16188 (n_8179, n8650);
  and g16189 (n8651, n680, n_8179);
  not g16190 (n_8180, n8651);
  and g16191 (n8652, n684, n_8180);
  not g16192 (n_8181, n8652);
  and g16193 (n8653, n688, n_8181);
  not g16194 (n_8182, n8653);
  and g16195 (n8654, n692, n_8182);
  not g16196 (n_8183, n8654);
  and g16197 (n8655, n696, n_8183);
  not g16198 (n_8184, n8655);
  and g16199 (n8656, n700, n_8184);
  not g16200 (n_8185, n8656);
  and g16201 (n8657, n704, n_8185);
  not g16202 (n_8186, n8657);
  and g16203 (n8658, n708, n_8186);
  not g16204 (n_8187, n8658);
  and g16205 (n8659, n712, n_8187);
  not g16206 (n_8188, n8659);
  and g16207 (n8660, n716, n_8188);
  not g16208 (n_8189, n8660);
  and g16209 (n8661, n720, n_8189);
  not g16210 (n_8190, n8661);
  and g16211 (n8662, n1484, n_8190);
  not g16212 (n_8191, n8662);
  and g16213 (n8663, n1486, n_8191);
  not g16214 (n_8192, n8663);
  and g16215 (n8664, n1750, n_8192);
  not g16216 (n_8193, n8664);
  and g16217 (n8665, n731, n_8193);
  not g16218 (n_8194, n8665);
  and g16219 (n8666, n735, n_8194);
  not g16220 (n_8195, n8666);
  and g16221 (n8667, n739, n_8195);
  not g16222 (n_8196, n8667);
  and g16223 (n8668, n743, n_8196);
  not g16224 (n_8197, n8668);
  and g16225 (n8669, n747, n_8197);
  not g16226 (n_8198, n8669);
  and g16227 (n8670, n751, n_8198);
  not g16228 (n_8199, n8670);
  and g16229 (n8671, n755, n_8199);
  not g16230 (n_8200, n8671);
  and g16231 (n8672, n759, n_8200);
  not g16232 (n_8201, n8672);
  and g16233 (n8673, n763, n_8201);
  not g16234 (n_8202, n8673);
  and g16235 (n8674, n767, n_8202);
  not g16236 (n_8203, n8674);
  and g16237 (n8675, n771, n_8203);
  not g16238 (n_8204, n8675);
  and g16239 (n8676, n775, n_8204);
  not g16240 (n_8205, n8676);
  and g16241 (n8677, n779, n_8205);
  not g16242 (n_8206, n8677);
  and g16243 (n8678, n783, n_8206);
  not g16244 (n_8207, n8678);
  and g16245 (n8679, n787, n_8207);
  not g16246 (n_8208, n8679);
  and g16247 (n8680, n791, n_8208);
  not g16248 (n_8209, n8680);
  and g16249 (n8681, n795, n_8209);
  not g16250 (n_8210, n8681);
  and g16251 (n8682, n799, n_8210);
  not g16252 (n_8211, n8682);
  and g16253 (n8683, n803, n_8211);
  not g16254 (n_8212, n8683);
  and g16255 (n8684, n807, n_8212);
  not g16256 (n_8213, n8684);
  and g16257 (n8685, n811, n_8213);
  not g16258 (n_8214, n8685);
  and g16259 (n8686, n815, n_8214);
  not g16260 (n_8215, n8686);
  and g16261 (n8687, n819, n_8215);
  not g16262 (n_8216, n8687);
  and g16263 (n8688, n823, n_8216);
  not g16264 (n_8217, n8688);
  and g16265 (n8689, n827, n_8217);
  not g16266 (n_8218, n8689);
  and g16267 (n8690, n831, n_8218);
  not g16268 (n_8219, n8690);
  and g16269 (n8691, n835, n_8219);
  not g16270 (n_8220, n8691);
  and g16271 (n8692, n839, n_8220);
  not g16272 (n_8221, n8692);
  and g16273 (n8693, n843, n_8221);
  not g16274 (n_8222, n8693);
  and g16275 (n8694, n847, n_8222);
  not g16276 (n_8223, n8694);
  and g16277 (n8695, n851, n_8223);
  not g16278 (n_8224, n8695);
  and g16279 (n8696, n855, n_8224);
  not g16280 (n_8225, n8696);
  and g16281 (n8697, n859, n_8225);
  not g16282 (n_8226, n8697);
  and g16283 (n8698, n863, n_8226);
  not g16284 (n_8227, n8698);
  and g16285 (n8699, n867, n_8227);
  not g16286 (n_8228, n8699);
  and g16287 (n8700, n871, n_8228);
  not g16288 (n_8229, n8700);
  and g16289 (n8701, n875, n_8229);
  not g16290 (n_8230, n8701);
  and g16291 (n8702, n879, n_8230);
  not g16292 (n_8231, n8702);
  and g16293 (n8703, n883, n_8231);
  not g16294 (n_8232, n8703);
  and g16295 (n8704, n887, n_8232);
  not g16296 (n_8233, n8704);
  and g16297 (n8705, n891, n_8233);
  not g16298 (n_8234, n8705);
  and g16299 (n8706, n895, n_8234);
  not g16300 (n_8235, n8706);
  and g16301 (n8707, n899, n_8235);
  not g16302 (n_8236, n8707);
  and g16303 (n8708, n903, n_8236);
  not g16304 (n_8237, n8708);
  and g16305 (n8709, n907, n_8237);
  not g16306 (n_8238, n8709);
  and g16307 (n8710, n911, n_8238);
  not g16308 (n_8239, n8710);
  and g16309 (n8711, n915, n_8239);
  not g16310 (n_8240, n8711);
  and g16311 (n8712, n919, n_8240);
  not g16312 (n_8241, n8712);
  and g16313 (n8713, n923, n_8241);
  not g16314 (n_8242, n8713);
  and g16315 (n8714, n927, n_8242);
  not g16316 (n_8243, n8714);
  and g16317 (n8715, n931, n_8243);
  not g16318 (n_8244, n8715);
  and g16319 (n8716, n935, n_8244);
  not g16320 (n_8245, n8716);
  and g16321 (n8717, n939, n_8245);
  not g16322 (n_8246, n8717);
  and g16323 (n8718, n943, n_8246);
  not g16324 (n_8247, n8718);
  and g16325 (n8719, n947, n_8247);
  and g16326 (n8720, \req[87] , n_767);
  not g16327 (n_8248, n8719);
  and g16328 (\grant[87] , n_8248, n8720);
  not g16329 (n_8249, n1291);
  and g16330 (n8722, n958, n_8249);
  not g16331 (n_8250, n8722);
  and g16332 (n8723, n963, n_8250);
  not g16333 (n_8251, n8723);
  and g16334 (n8724, n967, n_8251);
  not g16335 (n_8252, n8724);
  and g16336 (n8725, n971, n_8252);
  not g16337 (n_8253, n8725);
  and g16338 (n8726, n975, n_8253);
  not g16339 (n_8254, n8726);
  and g16340 (n8727, n979, n_8254);
  not g16341 (n_8255, n8727);
  and g16342 (n8728, n983, n_8255);
  not g16343 (n_8256, n8728);
  and g16344 (n8729, n987, n_8256);
  not g16345 (n_8257, n8729);
  and g16346 (n8730, n991, n_8257);
  not g16347 (n_8258, n8730);
  and g16348 (n8731, n995, n_8258);
  not g16349 (n_8259, n8731);
  and g16350 (n8732, n999, n_8259);
  not g16351 (n_8260, n8732);
  and g16352 (n8733, n1003, n_8260);
  not g16353 (n_8261, n8733);
  and g16354 (n8734, n1007, n_8261);
  not g16355 (n_8262, n8734);
  and g16356 (n8735, n1011, n_8262);
  not g16357 (n_8263, n8735);
  and g16358 (n8736, n1015, n_8263);
  not g16359 (n_8264, n8736);
  and g16360 (n8737, n1019, n_8264);
  not g16361 (n_8265, n8737);
  and g16362 (n8738, n1023, n_8265);
  not g16363 (n_8266, n8738);
  and g16364 (n8739, n1027, n_8266);
  not g16365 (n_8267, n8739);
  and g16366 (n8740, n1031, n_8267);
  not g16367 (n_8268, n8740);
  and g16368 (n8741, n1035, n_8268);
  not g16369 (n_8269, n8741);
  and g16370 (n8742, n1039, n_8269);
  not g16371 (n_8270, n8742);
  and g16372 (n8743, n1043, n_8270);
  not g16373 (n_8271, n8743);
  and g16374 (n8744, n1047, n_8271);
  not g16375 (n_8272, n8744);
  and g16376 (n8745, n1051, n_8272);
  not g16377 (n_8273, n8745);
  and g16378 (n8746, n1055, n_8273);
  not g16379 (n_8274, n8746);
  and g16380 (n8747, n1059, n_8274);
  not g16381 (n_8275, n8747);
  and g16382 (n8748, n1574, n_8275);
  not g16383 (n_8276, n8748);
  and g16384 (n8749, n1576, n_8276);
  not g16385 (n_8277, n8749);
  and g16386 (n8750, n1837, n_8277);
  not g16387 (n_8278, n8750);
  and g16388 (n8751, n1068, n_8278);
  not g16389 (n_8279, n8751);
  and g16390 (n8752, n1072, n_8279);
  not g16391 (n_8280, n8752);
  and g16392 (n8753, n1076, n_8280);
  not g16393 (n_8281, n8753);
  and g16394 (n8754, n1080, n_8281);
  not g16395 (n_8282, n8754);
  and g16396 (n8755, n1084, n_8282);
  not g16397 (n_8283, n8755);
  and g16398 (n8756, n1088, n_8283);
  not g16399 (n_8284, n8756);
  and g16400 (n8757, n1092, n_8284);
  not g16401 (n_8285, n8757);
  and g16402 (n8758, n1096, n_8285);
  not g16403 (n_8286, n8758);
  and g16404 (n8759, n1100, n_8286);
  not g16405 (n_8287, n8759);
  and g16406 (n8760, n1104, n_8287);
  not g16407 (n_8288, n8760);
  and g16408 (n8761, n1108, n_8288);
  not g16409 (n_8289, n8761);
  and g16410 (n8762, n1112, n_8289);
  not g16411 (n_8290, n8762);
  and g16412 (n8763, n1116, n_8290);
  not g16413 (n_8291, n8763);
  and g16414 (n8764, n1120, n_8291);
  not g16415 (n_8292, n8764);
  and g16416 (n8765, n1124, n_8292);
  not g16417 (n_8293, n8765);
  and g16418 (n8766, n1128, n_8293);
  not g16419 (n_8294, n8766);
  and g16420 (n8767, n1132, n_8294);
  not g16421 (n_8295, n8767);
  and g16422 (n8768, n1136, n_8295);
  not g16423 (n_8296, n8768);
  and g16424 (n8769, n1140, n_8296);
  not g16425 (n_8297, n8769);
  and g16426 (n8770, n1144, n_8297);
  not g16427 (n_8298, n8770);
  and g16428 (n8771, n1148, n_8298);
  not g16429 (n_8299, n8771);
  and g16430 (n8772, n1152, n_8299);
  not g16431 (n_8300, n8772);
  and g16432 (n8773, n1156, n_8300);
  not g16433 (n_8301, n8773);
  and g16434 (n8774, n1160, n_8301);
  not g16435 (n_8302, n8774);
  and g16436 (n8775, n1164, n_8302);
  not g16437 (n_8303, n8775);
  and g16438 (n8776, n1168, n_8303);
  not g16439 (n_8304, n8776);
  and g16440 (n8777, n1172, n_8304);
  not g16441 (n_8305, n8777);
  and g16442 (n8778, n1176, n_8305);
  not g16443 (n_8306, n8778);
  and g16444 (n8779, n1180, n_8306);
  not g16445 (n_8307, n8779);
  and g16446 (n8780, n1184, n_8307);
  not g16447 (n_8308, n8780);
  and g16448 (n8781, n1188, n_8308);
  not g16449 (n_8309, n8781);
  and g16450 (n8782, n1192, n_8309);
  not g16451 (n_8310, n8782);
  and g16452 (n8783, n1196, n_8310);
  not g16453 (n_8311, n8783);
  and g16454 (n8784, n1200, n_8311);
  not g16455 (n_8312, n8784);
  and g16456 (n8785, n1204, n_8312);
  not g16457 (n_8313, n8785);
  and g16458 (n8786, n1208, n_8313);
  not g16459 (n_8314, n8786);
  and g16460 (n8787, n1212, n_8314);
  not g16461 (n_8315, n8787);
  and g16462 (n8788, n1216, n_8315);
  not g16463 (n_8316, n8788);
  and g16464 (n8789, n1220, n_8316);
  not g16465 (n_8317, n8789);
  and g16466 (n8790, n1224, n_8317);
  not g16467 (n_8318, n8790);
  and g16468 (n8791, n1228, n_8318);
  not g16469 (n_8319, n8791);
  and g16470 (n8792, n1232, n_8319);
  not g16471 (n_8320, n8792);
  and g16472 (n8793, n1236, n_8320);
  not g16473 (n_8321, n8793);
  and g16474 (n8794, n1240, n_8321);
  not g16475 (n_8322, n8794);
  and g16476 (n8795, n1244, n_8322);
  not g16477 (n_8323, n8795);
  and g16478 (n8796, n1248, n_8323);
  not g16479 (n_8324, n8796);
  and g16480 (n8797, n1252, n_8324);
  not g16481 (n_8325, n8797);
  and g16482 (n8798, n1256, n_8325);
  not g16483 (n_8326, n8798);
  and g16484 (n8799, n1260, n_8326);
  not g16485 (n_8327, n8799);
  and g16486 (n8800, n1264, n_8327);
  not g16487 (n_8328, n8800);
  and g16488 (n8801, n1268, n_8328);
  not g16489 (n_8329, n8801);
  and g16490 (n8802, n1272, n_8329);
  not g16491 (n_8330, n8802);
  and g16492 (n8803, n1276, n_8330);
  not g16493 (n_8331, n8803);
  and g16494 (n8804, n1280, n_8331);
  not g16495 (n_8332, n8804);
  and g16496 (n8805, n1284, n_8332);
  and g16497 (n8806, \req[88] , n_963);
  not g16498 (n_8333, n8805);
  and g16499 (\grant[88] , n_8333, n8806);
  not g16500 (n_8334, n623);
  and g16501 (n8808, n_8334, n1295);
  not g16502 (n_8335, n8808);
  and g16503 (n8809, n1300, n_8335);
  not g16504 (n_8336, n8809);
  and g16505 (n8810, n1304, n_8336);
  not g16506 (n_8337, n8810);
  and g16507 (n8811, n1308, n_8337);
  not g16508 (n_8338, n8811);
  and g16509 (n8812, n1312, n_8338);
  not g16510 (n_8339, n8812);
  and g16511 (n8813, n1316, n_8339);
  not g16512 (n_8340, n8813);
  and g16513 (n8814, n1320, n_8340);
  not g16514 (n_8341, n8814);
  and g16515 (n8815, n1324, n_8341);
  not g16516 (n_8342, n8815);
  and g16517 (n8816, n1328, n_8342);
  not g16518 (n_8343, n8816);
  and g16519 (n8817, n1332, n_8343);
  not g16520 (n_8344, n8817);
  and g16521 (n8818, n1336, n_8344);
  not g16522 (n_8345, n8818);
  and g16523 (n8819, n1340, n_8345);
  not g16524 (n_8346, n8819);
  and g16525 (n8820, n1344, n_8346);
  not g16526 (n_8347, n8820);
  and g16527 (n8821, n1348, n_8347);
  not g16528 (n_8348, n8821);
  and g16529 (n8822, n1352, n_8348);
  not g16530 (n_8349, n8822);
  and g16531 (n8823, n1356, n_8349);
  not g16532 (n_8350, n8823);
  and g16533 (n8824, n1360, n_8350);
  not g16534 (n_8351, n8824);
  and g16535 (n8825, n1364, n_8351);
  not g16536 (n_8352, n8825);
  and g16537 (n8826, n1368, n_8352);
  not g16538 (n_8353, n8826);
  and g16539 (n8827, n1372, n_8353);
  not g16540 (n_8354, n8827);
  and g16541 (n8828, n1376, n_8354);
  not g16542 (n_8355, n8828);
  and g16543 (n8829, n1380, n_8355);
  not g16544 (n_8356, n8829);
  and g16545 (n8830, n1384, n_8356);
  not g16546 (n_8357, n8830);
  and g16547 (n8831, n1388, n_8357);
  not g16548 (n_8358, n8831);
  and g16549 (n8832, n1392, n_8358);
  not g16550 (n_8359, n8832);
  and g16551 (n8833, n1396, n_8359);
  not g16552 (n_8360, n8833);
  and g16553 (n8834, n1663, n_8360);
  not g16554 (n_8361, n8834);
  and g16555 (n8835, n392, n_8361);
  not g16556 (n_8362, n8835);
  and g16557 (n8836, n396, n_8362);
  not g16558 (n_8363, n8836);
  and g16559 (n8837, n400, n_8363);
  not g16560 (n_8364, n8837);
  and g16561 (n8838, n404, n_8364);
  not g16562 (n_8365, n8838);
  and g16563 (n8839, n408, n_8365);
  not g16564 (n_8366, n8839);
  and g16565 (n8840, n412, n_8366);
  not g16566 (n_8367, n8840);
  and g16567 (n8841, n416, n_8367);
  not g16568 (n_8368, n8841);
  and g16569 (n8842, n420, n_8368);
  not g16570 (n_8369, n8842);
  and g16571 (n8843, n424, n_8369);
  not g16572 (n_8370, n8843);
  and g16573 (n8844, n428, n_8370);
  not g16574 (n_8371, n8844);
  and g16575 (n8845, n432, n_8371);
  not g16576 (n_8372, n8845);
  and g16577 (n8846, n436, n_8372);
  not g16578 (n_8373, n8846);
  and g16579 (n8847, n440, n_8373);
  not g16580 (n_8374, n8847);
  and g16581 (n8848, n444, n_8374);
  not g16582 (n_8375, n8848);
  and g16583 (n8849, n448, n_8375);
  not g16584 (n_8376, n8849);
  and g16585 (n8850, n452, n_8376);
  not g16586 (n_8377, n8850);
  and g16587 (n8851, n456, n_8377);
  not g16588 (n_8378, n8851);
  and g16589 (n8852, n460, n_8378);
  not g16590 (n_8379, n8852);
  and g16591 (n8853, n464, n_8379);
  not g16592 (n_8380, n8853);
  and g16593 (n8854, n468, n_8380);
  not g16594 (n_8381, n8854);
  and g16595 (n8855, n472, n_8381);
  not g16596 (n_8382, n8855);
  and g16597 (n8856, n476, n_8382);
  not g16598 (n_8383, n8856);
  and g16599 (n8857, n480, n_8383);
  not g16600 (n_8384, n8857);
  and g16601 (n8858, n484, n_8384);
  not g16602 (n_8385, n8858);
  and g16603 (n8859, n488, n_8385);
  not g16604 (n_8386, n8859);
  and g16605 (n8860, n492, n_8386);
  not g16606 (n_8387, n8860);
  and g16607 (n8861, n496, n_8387);
  not g16608 (n_8388, n8861);
  and g16609 (n8862, n500, n_8388);
  not g16610 (n_8389, n8862);
  and g16611 (n8863, n504, n_8389);
  not g16612 (n_8390, n8863);
  and g16613 (n8864, n508, n_8390);
  not g16614 (n_8391, n8864);
  and g16615 (n8865, n512, n_8391);
  not g16616 (n_8392, n8865);
  and g16617 (n8866, n516, n_8392);
  not g16618 (n_8393, n8866);
  and g16619 (n8867, n520, n_8393);
  not g16620 (n_8394, n8867);
  and g16621 (n8868, n524, n_8394);
  not g16622 (n_8395, n8868);
  and g16623 (n8869, n528, n_8395);
  not g16624 (n_8396, n8869);
  and g16625 (n8870, n532, n_8396);
  not g16626 (n_8397, n8870);
  and g16627 (n8871, n536, n_8397);
  not g16628 (n_8398, n8871);
  and g16629 (n8872, n540, n_8398);
  not g16630 (n_8399, n8872);
  and g16631 (n8873, n544, n_8399);
  not g16632 (n_8400, n8873);
  and g16633 (n8874, n548, n_8400);
  not g16634 (n_8401, n8874);
  and g16635 (n8875, n552, n_8401);
  not g16636 (n_8402, n8875);
  and g16637 (n8876, n556, n_8402);
  not g16638 (n_8403, n8876);
  and g16639 (n8877, n560, n_8403);
  not g16640 (n_8404, n8877);
  and g16641 (n8878, n564, n_8404);
  not g16642 (n_8405, n8878);
  and g16643 (n8879, n568, n_8405);
  not g16644 (n_8406, n8879);
  and g16645 (n8880, n572, n_8406);
  not g16646 (n_8407, n8880);
  and g16647 (n8881, n576, n_8407);
  not g16648 (n_8408, n8881);
  and g16649 (n8882, n580, n_8408);
  not g16650 (n_8409, n8882);
  and g16651 (n8883, n584, n_8409);
  not g16652 (n_8410, n8883);
  and g16653 (n8884, n588, n_8410);
  not g16654 (n_8411, n8884);
  and g16655 (n8885, n592, n_8411);
  not g16656 (n_8412, n8885);
  and g16657 (n8886, n596, n_8412);
  not g16658 (n_8413, n8886);
  and g16659 (n8887, n600, n_8413);
  not g16660 (n_8414, n8887);
  and g16661 (n8888, n604, n_8414);
  not g16662 (n_8415, n8888);
  and g16663 (n8889, n608, n_8415);
  not g16664 (n_8416, n8889);
  and g16665 (n8890, n612, n_8416);
  not g16666 (n_8417, n8890);
  and g16667 (n8891, n616, n_8417);
  and g16668 (n8892, \req[89] , n_416);
  not g16669 (n_8418, n8891);
  and g16670 (\grant[89] , n_8418, n8892);
  not g16671 (n_8419, n962);
  and g16672 (n8894, n627, n_8419);
  not g16673 (n_8420, n8894);
  and g16674 (n8895, n632, n_8420);
  not g16675 (n_8421, n8895);
  and g16676 (n8896, n636, n_8421);
  not g16677 (n_8422, n8896);
  and g16678 (n8897, n640, n_8422);
  not g16679 (n_8423, n8897);
  and g16680 (n8898, n644, n_8423);
  not g16681 (n_8424, n8898);
  and g16682 (n8899, n648, n_8424);
  not g16683 (n_8425, n8899);
  and g16684 (n8900, n652, n_8425);
  not g16685 (n_8426, n8900);
  and g16686 (n8901, n656, n_8426);
  not g16687 (n_8427, n8901);
  and g16688 (n8902, n660, n_8427);
  not g16689 (n_8428, n8902);
  and g16690 (n8903, n664, n_8428);
  not g16691 (n_8429, n8903);
  and g16692 (n8904, n668, n_8429);
  not g16693 (n_8430, n8904);
  and g16694 (n8905, n672, n_8430);
  not g16695 (n_8431, n8905);
  and g16696 (n8906, n676, n_8431);
  not g16697 (n_8432, n8906);
  and g16698 (n8907, n680, n_8432);
  not g16699 (n_8433, n8907);
  and g16700 (n8908, n684, n_8433);
  not g16701 (n_8434, n8908);
  and g16702 (n8909, n688, n_8434);
  not g16703 (n_8435, n8909);
  and g16704 (n8910, n692, n_8435);
  not g16705 (n_8436, n8910);
  and g16706 (n8911, n696, n_8436);
  not g16707 (n_8437, n8911);
  and g16708 (n8912, n700, n_8437);
  not g16709 (n_8438, n8912);
  and g16710 (n8913, n704, n_8438);
  not g16711 (n_8439, n8913);
  and g16712 (n8914, n708, n_8439);
  not g16713 (n_8440, n8914);
  and g16714 (n8915, n712, n_8440);
  not g16715 (n_8441, n8915);
  and g16716 (n8916, n716, n_8441);
  not g16717 (n_8442, n8916);
  and g16718 (n8917, n720, n_8442);
  not g16719 (n_8443, n8917);
  and g16720 (n8918, n1484, n_8443);
  not g16721 (n_8444, n8918);
  and g16722 (n8919, n1486, n_8444);
  not g16723 (n_8445, n8919);
  and g16724 (n8920, n1750, n_8445);
  not g16725 (n_8446, n8920);
  and g16726 (n8921, n731, n_8446);
  not g16727 (n_8447, n8921);
  and g16728 (n8922, n735, n_8447);
  not g16729 (n_8448, n8922);
  and g16730 (n8923, n739, n_8448);
  not g16731 (n_8449, n8923);
  and g16732 (n8924, n743, n_8449);
  not g16733 (n_8450, n8924);
  and g16734 (n8925, n747, n_8450);
  not g16735 (n_8451, n8925);
  and g16736 (n8926, n751, n_8451);
  not g16737 (n_8452, n8926);
  and g16738 (n8927, n755, n_8452);
  not g16739 (n_8453, n8927);
  and g16740 (n8928, n759, n_8453);
  not g16741 (n_8454, n8928);
  and g16742 (n8929, n763, n_8454);
  not g16743 (n_8455, n8929);
  and g16744 (n8930, n767, n_8455);
  not g16745 (n_8456, n8930);
  and g16746 (n8931, n771, n_8456);
  not g16747 (n_8457, n8931);
  and g16748 (n8932, n775, n_8457);
  not g16749 (n_8458, n8932);
  and g16750 (n8933, n779, n_8458);
  not g16751 (n_8459, n8933);
  and g16752 (n8934, n783, n_8459);
  not g16753 (n_8460, n8934);
  and g16754 (n8935, n787, n_8460);
  not g16755 (n_8461, n8935);
  and g16756 (n8936, n791, n_8461);
  not g16757 (n_8462, n8936);
  and g16758 (n8937, n795, n_8462);
  not g16759 (n_8463, n8937);
  and g16760 (n8938, n799, n_8463);
  not g16761 (n_8464, n8938);
  and g16762 (n8939, n803, n_8464);
  not g16763 (n_8465, n8939);
  and g16764 (n8940, n807, n_8465);
  not g16765 (n_8466, n8940);
  and g16766 (n8941, n811, n_8466);
  not g16767 (n_8467, n8941);
  and g16768 (n8942, n815, n_8467);
  not g16769 (n_8468, n8942);
  and g16770 (n8943, n819, n_8468);
  not g16771 (n_8469, n8943);
  and g16772 (n8944, n823, n_8469);
  not g16773 (n_8470, n8944);
  and g16774 (n8945, n827, n_8470);
  not g16775 (n_8471, n8945);
  and g16776 (n8946, n831, n_8471);
  not g16777 (n_8472, n8946);
  and g16778 (n8947, n835, n_8472);
  not g16779 (n_8473, n8947);
  and g16780 (n8948, n839, n_8473);
  not g16781 (n_8474, n8948);
  and g16782 (n8949, n843, n_8474);
  not g16783 (n_8475, n8949);
  and g16784 (n8950, n847, n_8475);
  not g16785 (n_8476, n8950);
  and g16786 (n8951, n851, n_8476);
  not g16787 (n_8477, n8951);
  and g16788 (n8952, n855, n_8477);
  not g16789 (n_8478, n8952);
  and g16790 (n8953, n859, n_8478);
  not g16791 (n_8479, n8953);
  and g16792 (n8954, n863, n_8479);
  not g16793 (n_8480, n8954);
  and g16794 (n8955, n867, n_8480);
  not g16795 (n_8481, n8955);
  and g16796 (n8956, n871, n_8481);
  not g16797 (n_8482, n8956);
  and g16798 (n8957, n875, n_8482);
  not g16799 (n_8483, n8957);
  and g16800 (n8958, n879, n_8483);
  not g16801 (n_8484, n8958);
  and g16802 (n8959, n883, n_8484);
  not g16803 (n_8485, n8959);
  and g16804 (n8960, n887, n_8485);
  not g16805 (n_8486, n8960);
  and g16806 (n8961, n891, n_8486);
  not g16807 (n_8487, n8961);
  and g16808 (n8962, n895, n_8487);
  not g16809 (n_8488, n8962);
  and g16810 (n8963, n899, n_8488);
  not g16811 (n_8489, n8963);
  and g16812 (n8964, n903, n_8489);
  not g16813 (n_8490, n8964);
  and g16814 (n8965, n907, n_8490);
  not g16815 (n_8491, n8965);
  and g16816 (n8966, n911, n_8491);
  not g16817 (n_8492, n8966);
  and g16818 (n8967, n915, n_8492);
  not g16819 (n_8493, n8967);
  and g16820 (n8968, n919, n_8493);
  not g16821 (n_8494, n8968);
  and g16822 (n8969, n923, n_8494);
  not g16823 (n_8495, n8969);
  and g16824 (n8970, n927, n_8495);
  not g16825 (n_8496, n8970);
  and g16826 (n8971, n931, n_8496);
  not g16827 (n_8497, n8971);
  and g16828 (n8972, n935, n_8497);
  not g16829 (n_8498, n8972);
  and g16830 (n8973, n939, n_8498);
  not g16831 (n_8499, n8973);
  and g16832 (n8974, n943, n_8499);
  not g16833 (n_8500, n8974);
  and g16834 (n8975, n947, n_8500);
  not g16835 (n_8501, n8975);
  and g16836 (n8976, n951, n_8501);
  not g16837 (n_8502, n8976);
  and g16838 (n8977, n955, n_8502);
  and g16839 (n8978, \req[90] , n_773);
  not g16840 (n_8503, n8977);
  and g16841 (\grant[90] , n_8503, n8978);
  not g16842 (n_8504, n1299);
  and g16843 (n8980, n966, n_8504);
  not g16844 (n_8505, n8980);
  and g16845 (n8981, n971, n_8505);
  not g16846 (n_8506, n8981);
  and g16847 (n8982, n975, n_8506);
  not g16848 (n_8507, n8982);
  and g16849 (n8983, n979, n_8507);
  not g16850 (n_8508, n8983);
  and g16851 (n8984, n983, n_8508);
  not g16852 (n_8509, n8984);
  and g16853 (n8985, n987, n_8509);
  not g16854 (n_8510, n8985);
  and g16855 (n8986, n991, n_8510);
  not g16856 (n_8511, n8986);
  and g16857 (n8987, n995, n_8511);
  not g16858 (n_8512, n8987);
  and g16859 (n8988, n999, n_8512);
  not g16860 (n_8513, n8988);
  and g16861 (n8989, n1003, n_8513);
  not g16862 (n_8514, n8989);
  and g16863 (n8990, n1007, n_8514);
  not g16864 (n_8515, n8990);
  and g16865 (n8991, n1011, n_8515);
  not g16866 (n_8516, n8991);
  and g16867 (n8992, n1015, n_8516);
  not g16868 (n_8517, n8992);
  and g16869 (n8993, n1019, n_8517);
  not g16870 (n_8518, n8993);
  and g16871 (n8994, n1023, n_8518);
  not g16872 (n_8519, n8994);
  and g16873 (n8995, n1027, n_8519);
  not g16874 (n_8520, n8995);
  and g16875 (n8996, n1031, n_8520);
  not g16876 (n_8521, n8996);
  and g16877 (n8997, n1035, n_8521);
  not g16878 (n_8522, n8997);
  and g16879 (n8998, n1039, n_8522);
  not g16880 (n_8523, n8998);
  and g16881 (n8999, n1043, n_8523);
  not g16882 (n_8524, n8999);
  and g16883 (n9000, n1047, n_8524);
  not g16884 (n_8525, n9000);
  and g16885 (n9001, n1051, n_8525);
  not g16886 (n_8526, n9001);
  and g16887 (n9002, n1055, n_8526);
  not g16888 (n_8527, n9002);
  and g16889 (n9003, n1059, n_8527);
  not g16890 (n_8528, n9003);
  and g16891 (n9004, n1574, n_8528);
  not g16892 (n_8529, n9004);
  and g16893 (n9005, n1576, n_8529);
  not g16894 (n_8530, n9005);
  and g16895 (n9006, n1837, n_8530);
  not g16896 (n_8531, n9006);
  and g16897 (n9007, n1068, n_8531);
  not g16898 (n_8532, n9007);
  and g16899 (n9008, n1072, n_8532);
  not g16900 (n_8533, n9008);
  and g16901 (n9009, n1076, n_8533);
  not g16902 (n_8534, n9009);
  and g16903 (n9010, n1080, n_8534);
  not g16904 (n_8535, n9010);
  and g16905 (n9011, n1084, n_8535);
  not g16906 (n_8536, n9011);
  and g16907 (n9012, n1088, n_8536);
  not g16908 (n_8537, n9012);
  and g16909 (n9013, n1092, n_8537);
  not g16910 (n_8538, n9013);
  and g16911 (n9014, n1096, n_8538);
  not g16912 (n_8539, n9014);
  and g16913 (n9015, n1100, n_8539);
  not g16914 (n_8540, n9015);
  and g16915 (n9016, n1104, n_8540);
  not g16916 (n_8541, n9016);
  and g16917 (n9017, n1108, n_8541);
  not g16918 (n_8542, n9017);
  and g16919 (n9018, n1112, n_8542);
  not g16920 (n_8543, n9018);
  and g16921 (n9019, n1116, n_8543);
  not g16922 (n_8544, n9019);
  and g16923 (n9020, n1120, n_8544);
  not g16924 (n_8545, n9020);
  and g16925 (n9021, n1124, n_8545);
  not g16926 (n_8546, n9021);
  and g16927 (n9022, n1128, n_8546);
  not g16928 (n_8547, n9022);
  and g16929 (n9023, n1132, n_8547);
  not g16930 (n_8548, n9023);
  and g16931 (n9024, n1136, n_8548);
  not g16932 (n_8549, n9024);
  and g16933 (n9025, n1140, n_8549);
  not g16934 (n_8550, n9025);
  and g16935 (n9026, n1144, n_8550);
  not g16936 (n_8551, n9026);
  and g16937 (n9027, n1148, n_8551);
  not g16938 (n_8552, n9027);
  and g16939 (n9028, n1152, n_8552);
  not g16940 (n_8553, n9028);
  and g16941 (n9029, n1156, n_8553);
  not g16942 (n_8554, n9029);
  and g16943 (n9030, n1160, n_8554);
  not g16944 (n_8555, n9030);
  and g16945 (n9031, n1164, n_8555);
  not g16946 (n_8556, n9031);
  and g16947 (n9032, n1168, n_8556);
  not g16948 (n_8557, n9032);
  and g16949 (n9033, n1172, n_8557);
  not g16950 (n_8558, n9033);
  and g16951 (n9034, n1176, n_8558);
  not g16952 (n_8559, n9034);
  and g16953 (n9035, n1180, n_8559);
  not g16954 (n_8560, n9035);
  and g16955 (n9036, n1184, n_8560);
  not g16956 (n_8561, n9036);
  and g16957 (n9037, n1188, n_8561);
  not g16958 (n_8562, n9037);
  and g16959 (n9038, n1192, n_8562);
  not g16960 (n_8563, n9038);
  and g16961 (n9039, n1196, n_8563);
  not g16962 (n_8564, n9039);
  and g16963 (n9040, n1200, n_8564);
  not g16964 (n_8565, n9040);
  and g16965 (n9041, n1204, n_8565);
  not g16966 (n_8566, n9041);
  and g16967 (n9042, n1208, n_8566);
  not g16968 (n_8567, n9042);
  and g16969 (n9043, n1212, n_8567);
  not g16970 (n_8568, n9043);
  and g16971 (n9044, n1216, n_8568);
  not g16972 (n_8569, n9044);
  and g16973 (n9045, n1220, n_8569);
  not g16974 (n_8570, n9045);
  and g16975 (n9046, n1224, n_8570);
  not g16976 (n_8571, n9046);
  and g16977 (n9047, n1228, n_8571);
  not g16978 (n_8572, n9047);
  and g16979 (n9048, n1232, n_8572);
  not g16980 (n_8573, n9048);
  and g16981 (n9049, n1236, n_8573);
  not g16982 (n_8574, n9049);
  and g16983 (n9050, n1240, n_8574);
  not g16984 (n_8575, n9050);
  and g16985 (n9051, n1244, n_8575);
  not g16986 (n_8576, n9051);
  and g16987 (n9052, n1248, n_8576);
  not g16988 (n_8577, n9052);
  and g16989 (n9053, n1252, n_8577);
  not g16990 (n_8578, n9053);
  and g16991 (n9054, n1256, n_8578);
  not g16992 (n_8579, n9054);
  and g16993 (n9055, n1260, n_8579);
  not g16994 (n_8580, n9055);
  and g16995 (n9056, n1264, n_8580);
  not g16996 (n_8581, n9056);
  and g16997 (n9057, n1268, n_8581);
  not g16998 (n_8582, n9057);
  and g16999 (n9058, n1272, n_8582);
  not g17000 (n_8583, n9058);
  and g17001 (n9059, n1276, n_8583);
  not g17002 (n_8584, n9059);
  and g17003 (n9060, n1280, n_8584);
  not g17004 (n_8585, n9060);
  and g17005 (n9061, n1284, n_8585);
  not g17006 (n_8586, n9061);
  and g17007 (n9062, n1288, n_8586);
  not g17008 (n_8587, n9062);
  and g17009 (n9063, n1292, n_8587);
  and g17010 (n9064, \req[91] , n_967);
  not g17011 (n_8588, n9063);
  and g17012 (\grant[91] , n_8588, n9064);
  not g17013 (n_8589, n631);
  and g17014 (n9066, n_8589, n1303);
  not g17015 (n_8590, n9066);
  and g17016 (n9067, n1308, n_8590);
  not g17017 (n_8591, n9067);
  and g17018 (n9068, n1312, n_8591);
  not g17019 (n_8592, n9068);
  and g17020 (n9069, n1316, n_8592);
  not g17021 (n_8593, n9069);
  and g17022 (n9070, n1320, n_8593);
  not g17023 (n_8594, n9070);
  and g17024 (n9071, n1324, n_8594);
  not g17025 (n_8595, n9071);
  and g17026 (n9072, n1328, n_8595);
  not g17027 (n_8596, n9072);
  and g17028 (n9073, n1332, n_8596);
  not g17029 (n_8597, n9073);
  and g17030 (n9074, n1336, n_8597);
  not g17031 (n_8598, n9074);
  and g17032 (n9075, n1340, n_8598);
  not g17033 (n_8599, n9075);
  and g17034 (n9076, n1344, n_8599);
  not g17035 (n_8600, n9076);
  and g17036 (n9077, n1348, n_8600);
  not g17037 (n_8601, n9077);
  and g17038 (n9078, n1352, n_8601);
  not g17039 (n_8602, n9078);
  and g17040 (n9079, n1356, n_8602);
  not g17041 (n_8603, n9079);
  and g17042 (n9080, n1360, n_8603);
  not g17043 (n_8604, n9080);
  and g17044 (n9081, n1364, n_8604);
  not g17045 (n_8605, n9081);
  and g17046 (n9082, n1368, n_8605);
  not g17047 (n_8606, n9082);
  and g17048 (n9083, n1372, n_8606);
  not g17049 (n_8607, n9083);
  and g17050 (n9084, n1376, n_8607);
  not g17051 (n_8608, n9084);
  and g17052 (n9085, n1380, n_8608);
  not g17053 (n_8609, n9085);
  and g17054 (n9086, n1384, n_8609);
  not g17055 (n_8610, n9086);
  and g17056 (n9087, n1388, n_8610);
  not g17057 (n_8611, n9087);
  and g17058 (n9088, n1392, n_8611);
  not g17059 (n_8612, n9088);
  and g17060 (n9089, n1396, n_8612);
  not g17061 (n_8613, n9089);
  and g17062 (n9090, n1663, n_8613);
  not g17063 (n_8614, n9090);
  and g17064 (n9091, n392, n_8614);
  not g17065 (n_8615, n9091);
  and g17066 (n9092, n396, n_8615);
  not g17067 (n_8616, n9092);
  and g17068 (n9093, n400, n_8616);
  not g17069 (n_8617, n9093);
  and g17070 (n9094, n404, n_8617);
  not g17071 (n_8618, n9094);
  and g17072 (n9095, n408, n_8618);
  not g17073 (n_8619, n9095);
  and g17074 (n9096, n412, n_8619);
  not g17075 (n_8620, n9096);
  and g17076 (n9097, n416, n_8620);
  not g17077 (n_8621, n9097);
  and g17078 (n9098, n420, n_8621);
  not g17079 (n_8622, n9098);
  and g17080 (n9099, n424, n_8622);
  not g17081 (n_8623, n9099);
  and g17082 (n9100, n428, n_8623);
  not g17083 (n_8624, n9100);
  and g17084 (n9101, n432, n_8624);
  not g17085 (n_8625, n9101);
  and g17086 (n9102, n436, n_8625);
  not g17087 (n_8626, n9102);
  and g17088 (n9103, n440, n_8626);
  not g17089 (n_8627, n9103);
  and g17090 (n9104, n444, n_8627);
  not g17091 (n_8628, n9104);
  and g17092 (n9105, n448, n_8628);
  not g17093 (n_8629, n9105);
  and g17094 (n9106, n452, n_8629);
  not g17095 (n_8630, n9106);
  and g17096 (n9107, n456, n_8630);
  not g17097 (n_8631, n9107);
  and g17098 (n9108, n460, n_8631);
  not g17099 (n_8632, n9108);
  and g17100 (n9109, n464, n_8632);
  not g17101 (n_8633, n9109);
  and g17102 (n9110, n468, n_8633);
  not g17103 (n_8634, n9110);
  and g17104 (n9111, n472, n_8634);
  not g17105 (n_8635, n9111);
  and g17106 (n9112, n476, n_8635);
  not g17107 (n_8636, n9112);
  and g17108 (n9113, n480, n_8636);
  not g17109 (n_8637, n9113);
  and g17110 (n9114, n484, n_8637);
  not g17111 (n_8638, n9114);
  and g17112 (n9115, n488, n_8638);
  not g17113 (n_8639, n9115);
  and g17114 (n9116, n492, n_8639);
  not g17115 (n_8640, n9116);
  and g17116 (n9117, n496, n_8640);
  not g17117 (n_8641, n9117);
  and g17118 (n9118, n500, n_8641);
  not g17119 (n_8642, n9118);
  and g17120 (n9119, n504, n_8642);
  not g17121 (n_8643, n9119);
  and g17122 (n9120, n508, n_8643);
  not g17123 (n_8644, n9120);
  and g17124 (n9121, n512, n_8644);
  not g17125 (n_8645, n9121);
  and g17126 (n9122, n516, n_8645);
  not g17127 (n_8646, n9122);
  and g17128 (n9123, n520, n_8646);
  not g17129 (n_8647, n9123);
  and g17130 (n9124, n524, n_8647);
  not g17131 (n_8648, n9124);
  and g17132 (n9125, n528, n_8648);
  not g17133 (n_8649, n9125);
  and g17134 (n9126, n532, n_8649);
  not g17135 (n_8650, n9126);
  and g17136 (n9127, n536, n_8650);
  not g17137 (n_8651, n9127);
  and g17138 (n9128, n540, n_8651);
  not g17139 (n_8652, n9128);
  and g17140 (n9129, n544, n_8652);
  not g17141 (n_8653, n9129);
  and g17142 (n9130, n548, n_8653);
  not g17143 (n_8654, n9130);
  and g17144 (n9131, n552, n_8654);
  not g17145 (n_8655, n9131);
  and g17146 (n9132, n556, n_8655);
  not g17147 (n_8656, n9132);
  and g17148 (n9133, n560, n_8656);
  not g17149 (n_8657, n9133);
  and g17150 (n9134, n564, n_8657);
  not g17151 (n_8658, n9134);
  and g17152 (n9135, n568, n_8658);
  not g17153 (n_8659, n9135);
  and g17154 (n9136, n572, n_8659);
  not g17155 (n_8660, n9136);
  and g17156 (n9137, n576, n_8660);
  not g17157 (n_8661, n9137);
  and g17158 (n9138, n580, n_8661);
  not g17159 (n_8662, n9138);
  and g17160 (n9139, n584, n_8662);
  not g17161 (n_8663, n9139);
  and g17162 (n9140, n588, n_8663);
  not g17163 (n_8664, n9140);
  and g17164 (n9141, n592, n_8664);
  not g17165 (n_8665, n9141);
  and g17166 (n9142, n596, n_8665);
  not g17167 (n_8666, n9142);
  and g17168 (n9143, n600, n_8666);
  not g17169 (n_8667, n9143);
  and g17170 (n9144, n604, n_8667);
  not g17171 (n_8668, n9144);
  and g17172 (n9145, n608, n_8668);
  not g17173 (n_8669, n9145);
  and g17174 (n9146, n612, n_8669);
  not g17175 (n_8670, n9146);
  and g17176 (n9147, n616, n_8670);
  not g17177 (n_8671, n9147);
  and g17178 (n9148, n620, n_8671);
  not g17179 (n_8672, n9148);
  and g17180 (n9149, n624, n_8672);
  and g17181 (n9150, \req[92] , n_430);
  not g17182 (n_8673, n9149);
  and g17183 (\grant[92] , n_8673, n9150);
  not g17184 (n_8674, n970);
  and g17185 (n9152, n635, n_8674);
  not g17186 (n_8675, n9152);
  and g17187 (n9153, n640, n_8675);
  not g17188 (n_8676, n9153);
  and g17189 (n9154, n644, n_8676);
  not g17190 (n_8677, n9154);
  and g17191 (n9155, n648, n_8677);
  not g17192 (n_8678, n9155);
  and g17193 (n9156, n652, n_8678);
  not g17194 (n_8679, n9156);
  and g17195 (n9157, n656, n_8679);
  not g17196 (n_8680, n9157);
  and g17197 (n9158, n660, n_8680);
  not g17198 (n_8681, n9158);
  and g17199 (n9159, n664, n_8681);
  not g17200 (n_8682, n9159);
  and g17201 (n9160, n668, n_8682);
  not g17202 (n_8683, n9160);
  and g17203 (n9161, n672, n_8683);
  not g17204 (n_8684, n9161);
  and g17205 (n9162, n676, n_8684);
  not g17206 (n_8685, n9162);
  and g17207 (n9163, n680, n_8685);
  not g17208 (n_8686, n9163);
  and g17209 (n9164, n684, n_8686);
  not g17210 (n_8687, n9164);
  and g17211 (n9165, n688, n_8687);
  not g17212 (n_8688, n9165);
  and g17213 (n9166, n692, n_8688);
  not g17214 (n_8689, n9166);
  and g17215 (n9167, n696, n_8689);
  not g17216 (n_8690, n9167);
  and g17217 (n9168, n700, n_8690);
  not g17218 (n_8691, n9168);
  and g17219 (n9169, n704, n_8691);
  not g17220 (n_8692, n9169);
  and g17221 (n9170, n708, n_8692);
  not g17222 (n_8693, n9170);
  and g17223 (n9171, n712, n_8693);
  not g17224 (n_8694, n9171);
  and g17225 (n9172, n716, n_8694);
  not g17226 (n_8695, n9172);
  and g17227 (n9173, n720, n_8695);
  not g17228 (n_8696, n9173);
  and g17229 (n9174, n1484, n_8696);
  not g17230 (n_8697, n9174);
  and g17231 (n9175, n1486, n_8697);
  not g17232 (n_8698, n9175);
  and g17233 (n9176, n1750, n_8698);
  not g17234 (n_8699, n9176);
  and g17235 (n9177, n731, n_8699);
  not g17236 (n_8700, n9177);
  and g17237 (n9178, n735, n_8700);
  not g17238 (n_8701, n9178);
  and g17239 (n9179, n739, n_8701);
  not g17240 (n_8702, n9179);
  and g17241 (n9180, n743, n_8702);
  not g17242 (n_8703, n9180);
  and g17243 (n9181, n747, n_8703);
  not g17244 (n_8704, n9181);
  and g17245 (n9182, n751, n_8704);
  not g17246 (n_8705, n9182);
  and g17247 (n9183, n755, n_8705);
  not g17248 (n_8706, n9183);
  and g17249 (n9184, n759, n_8706);
  not g17250 (n_8707, n9184);
  and g17251 (n9185, n763, n_8707);
  not g17252 (n_8708, n9185);
  and g17253 (n9186, n767, n_8708);
  not g17254 (n_8709, n9186);
  and g17255 (n9187, n771, n_8709);
  not g17256 (n_8710, n9187);
  and g17257 (n9188, n775, n_8710);
  not g17258 (n_8711, n9188);
  and g17259 (n9189, n779, n_8711);
  not g17260 (n_8712, n9189);
  and g17261 (n9190, n783, n_8712);
  not g17262 (n_8713, n9190);
  and g17263 (n9191, n787, n_8713);
  not g17264 (n_8714, n9191);
  and g17265 (n9192, n791, n_8714);
  not g17266 (n_8715, n9192);
  and g17267 (n9193, n795, n_8715);
  not g17268 (n_8716, n9193);
  and g17269 (n9194, n799, n_8716);
  not g17270 (n_8717, n9194);
  and g17271 (n9195, n803, n_8717);
  not g17272 (n_8718, n9195);
  and g17273 (n9196, n807, n_8718);
  not g17274 (n_8719, n9196);
  and g17275 (n9197, n811, n_8719);
  not g17276 (n_8720, n9197);
  and g17277 (n9198, n815, n_8720);
  not g17278 (n_8721, n9198);
  and g17279 (n9199, n819, n_8721);
  not g17280 (n_8722, n9199);
  and g17281 (n9200, n823, n_8722);
  not g17282 (n_8723, n9200);
  and g17283 (n9201, n827, n_8723);
  not g17284 (n_8724, n9201);
  and g17285 (n9202, n831, n_8724);
  not g17286 (n_8725, n9202);
  and g17287 (n9203, n835, n_8725);
  not g17288 (n_8726, n9203);
  and g17289 (n9204, n839, n_8726);
  not g17290 (n_8727, n9204);
  and g17291 (n9205, n843, n_8727);
  not g17292 (n_8728, n9205);
  and g17293 (n9206, n847, n_8728);
  not g17294 (n_8729, n9206);
  and g17295 (n9207, n851, n_8729);
  not g17296 (n_8730, n9207);
  and g17297 (n9208, n855, n_8730);
  not g17298 (n_8731, n9208);
  and g17299 (n9209, n859, n_8731);
  not g17300 (n_8732, n9209);
  and g17301 (n9210, n863, n_8732);
  not g17302 (n_8733, n9210);
  and g17303 (n9211, n867, n_8733);
  not g17304 (n_8734, n9211);
  and g17305 (n9212, n871, n_8734);
  not g17306 (n_8735, n9212);
  and g17307 (n9213, n875, n_8735);
  not g17308 (n_8736, n9213);
  and g17309 (n9214, n879, n_8736);
  not g17310 (n_8737, n9214);
  and g17311 (n9215, n883, n_8737);
  not g17312 (n_8738, n9215);
  and g17313 (n9216, n887, n_8738);
  not g17314 (n_8739, n9216);
  and g17315 (n9217, n891, n_8739);
  not g17316 (n_8740, n9217);
  and g17317 (n9218, n895, n_8740);
  not g17318 (n_8741, n9218);
  and g17319 (n9219, n899, n_8741);
  not g17320 (n_8742, n9219);
  and g17321 (n9220, n903, n_8742);
  not g17322 (n_8743, n9220);
  and g17323 (n9221, n907, n_8743);
  not g17324 (n_8744, n9221);
  and g17325 (n9222, n911, n_8744);
  not g17326 (n_8745, n9222);
  and g17327 (n9223, n915, n_8745);
  not g17328 (n_8746, n9223);
  and g17329 (n9224, n919, n_8746);
  not g17330 (n_8747, n9224);
  and g17331 (n9225, n923, n_8747);
  not g17332 (n_8748, n9225);
  and g17333 (n9226, n927, n_8748);
  not g17334 (n_8749, n9226);
  and g17335 (n9227, n931, n_8749);
  not g17336 (n_8750, n9227);
  and g17337 (n9228, n935, n_8750);
  not g17338 (n_8751, n9228);
  and g17339 (n9229, n939, n_8751);
  not g17340 (n_8752, n9229);
  and g17341 (n9230, n943, n_8752);
  not g17342 (n_8753, n9230);
  and g17343 (n9231, n947, n_8753);
  not g17344 (n_8754, n9231);
  and g17345 (n9232, n951, n_8754);
  not g17346 (n_8755, n9232);
  and g17347 (n9233, n955, n_8755);
  not g17348 (n_8756, n9233);
  and g17349 (n9234, n959, n_8756);
  not g17350 (n_8757, n9234);
  and g17351 (n9235, n963, n_8757);
  and g17352 (n9236, \req[93] , n_779);
  not g17353 (n_8758, n9235);
  and g17354 (\grant[93] , n_8758, n9236);
  not g17355 (n_8759, n1307);
  and g17356 (n9238, n974, n_8759);
  not g17357 (n_8760, n9238);
  and g17358 (n9239, n979, n_8760);
  not g17359 (n_8761, n9239);
  and g17360 (n9240, n983, n_8761);
  not g17361 (n_8762, n9240);
  and g17362 (n9241, n987, n_8762);
  not g17363 (n_8763, n9241);
  and g17364 (n9242, n991, n_8763);
  not g17365 (n_8764, n9242);
  and g17366 (n9243, n995, n_8764);
  not g17367 (n_8765, n9243);
  and g17368 (n9244, n999, n_8765);
  not g17369 (n_8766, n9244);
  and g17370 (n9245, n1003, n_8766);
  not g17371 (n_8767, n9245);
  and g17372 (n9246, n1007, n_8767);
  not g17373 (n_8768, n9246);
  and g17374 (n9247, n1011, n_8768);
  not g17375 (n_8769, n9247);
  and g17376 (n9248, n1015, n_8769);
  not g17377 (n_8770, n9248);
  and g17378 (n9249, n1019, n_8770);
  not g17379 (n_8771, n9249);
  and g17380 (n9250, n1023, n_8771);
  not g17381 (n_8772, n9250);
  and g17382 (n9251, n1027, n_8772);
  not g17383 (n_8773, n9251);
  and g17384 (n9252, n1031, n_8773);
  not g17385 (n_8774, n9252);
  and g17386 (n9253, n1035, n_8774);
  not g17387 (n_8775, n9253);
  and g17388 (n9254, n1039, n_8775);
  not g17389 (n_8776, n9254);
  and g17390 (n9255, n1043, n_8776);
  not g17391 (n_8777, n9255);
  and g17392 (n9256, n1047, n_8777);
  not g17393 (n_8778, n9256);
  and g17394 (n9257, n1051, n_8778);
  not g17395 (n_8779, n9257);
  and g17396 (n9258, n1055, n_8779);
  not g17397 (n_8780, n9258);
  and g17398 (n9259, n1059, n_8780);
  not g17399 (n_8781, n9259);
  and g17400 (n9260, n1574, n_8781);
  not g17401 (n_8782, n9260);
  and g17402 (n9261, n1576, n_8782);
  not g17403 (n_8783, n9261);
  and g17404 (n9262, n1837, n_8783);
  not g17405 (n_8784, n9262);
  and g17406 (n9263, n1068, n_8784);
  not g17407 (n_8785, n9263);
  and g17408 (n9264, n1072, n_8785);
  not g17409 (n_8786, n9264);
  and g17410 (n9265, n1076, n_8786);
  not g17411 (n_8787, n9265);
  and g17412 (n9266, n1080, n_8787);
  not g17413 (n_8788, n9266);
  and g17414 (n9267, n1084, n_8788);
  not g17415 (n_8789, n9267);
  and g17416 (n9268, n1088, n_8789);
  not g17417 (n_8790, n9268);
  and g17418 (n9269, n1092, n_8790);
  not g17419 (n_8791, n9269);
  and g17420 (n9270, n1096, n_8791);
  not g17421 (n_8792, n9270);
  and g17422 (n9271, n1100, n_8792);
  not g17423 (n_8793, n9271);
  and g17424 (n9272, n1104, n_8793);
  not g17425 (n_8794, n9272);
  and g17426 (n9273, n1108, n_8794);
  not g17427 (n_8795, n9273);
  and g17428 (n9274, n1112, n_8795);
  not g17429 (n_8796, n9274);
  and g17430 (n9275, n1116, n_8796);
  not g17431 (n_8797, n9275);
  and g17432 (n9276, n1120, n_8797);
  not g17433 (n_8798, n9276);
  and g17434 (n9277, n1124, n_8798);
  not g17435 (n_8799, n9277);
  and g17436 (n9278, n1128, n_8799);
  not g17437 (n_8800, n9278);
  and g17438 (n9279, n1132, n_8800);
  not g17439 (n_8801, n9279);
  and g17440 (n9280, n1136, n_8801);
  not g17441 (n_8802, n9280);
  and g17442 (n9281, n1140, n_8802);
  not g17443 (n_8803, n9281);
  and g17444 (n9282, n1144, n_8803);
  not g17445 (n_8804, n9282);
  and g17446 (n9283, n1148, n_8804);
  not g17447 (n_8805, n9283);
  and g17448 (n9284, n1152, n_8805);
  not g17449 (n_8806, n9284);
  and g17450 (n9285, n1156, n_8806);
  not g17451 (n_8807, n9285);
  and g17452 (n9286, n1160, n_8807);
  not g17453 (n_8808, n9286);
  and g17454 (n9287, n1164, n_8808);
  not g17455 (n_8809, n9287);
  and g17456 (n9288, n1168, n_8809);
  not g17457 (n_8810, n9288);
  and g17458 (n9289, n1172, n_8810);
  not g17459 (n_8811, n9289);
  and g17460 (n9290, n1176, n_8811);
  not g17461 (n_8812, n9290);
  and g17462 (n9291, n1180, n_8812);
  not g17463 (n_8813, n9291);
  and g17464 (n9292, n1184, n_8813);
  not g17465 (n_8814, n9292);
  and g17466 (n9293, n1188, n_8814);
  not g17467 (n_8815, n9293);
  and g17468 (n9294, n1192, n_8815);
  not g17469 (n_8816, n9294);
  and g17470 (n9295, n1196, n_8816);
  not g17471 (n_8817, n9295);
  and g17472 (n9296, n1200, n_8817);
  not g17473 (n_8818, n9296);
  and g17474 (n9297, n1204, n_8818);
  not g17475 (n_8819, n9297);
  and g17476 (n9298, n1208, n_8819);
  not g17477 (n_8820, n9298);
  and g17478 (n9299, n1212, n_8820);
  not g17479 (n_8821, n9299);
  and g17480 (n9300, n1216, n_8821);
  not g17481 (n_8822, n9300);
  and g17482 (n9301, n1220, n_8822);
  not g17483 (n_8823, n9301);
  and g17484 (n9302, n1224, n_8823);
  not g17485 (n_8824, n9302);
  and g17486 (n9303, n1228, n_8824);
  not g17487 (n_8825, n9303);
  and g17488 (n9304, n1232, n_8825);
  not g17489 (n_8826, n9304);
  and g17490 (n9305, n1236, n_8826);
  not g17491 (n_8827, n9305);
  and g17492 (n9306, n1240, n_8827);
  not g17493 (n_8828, n9306);
  and g17494 (n9307, n1244, n_8828);
  not g17495 (n_8829, n9307);
  and g17496 (n9308, n1248, n_8829);
  not g17497 (n_8830, n9308);
  and g17498 (n9309, n1252, n_8830);
  not g17499 (n_8831, n9309);
  and g17500 (n9310, n1256, n_8831);
  not g17501 (n_8832, n9310);
  and g17502 (n9311, n1260, n_8832);
  not g17503 (n_8833, n9311);
  and g17504 (n9312, n1264, n_8833);
  not g17505 (n_8834, n9312);
  and g17506 (n9313, n1268, n_8834);
  not g17507 (n_8835, n9313);
  and g17508 (n9314, n1272, n_8835);
  not g17509 (n_8836, n9314);
  and g17510 (n9315, n1276, n_8836);
  not g17511 (n_8837, n9315);
  and g17512 (n9316, n1280, n_8837);
  not g17513 (n_8838, n9316);
  and g17514 (n9317, n1284, n_8838);
  not g17515 (n_8839, n9317);
  and g17516 (n9318, n1288, n_8839);
  not g17517 (n_8840, n9318);
  and g17518 (n9319, n1292, n_8840);
  not g17519 (n_8841, n9319);
  and g17520 (n9320, n1296, n_8841);
  not g17521 (n_8842, n9320);
  and g17522 (n9321, n1300, n_8842);
  and g17523 (n9322, \req[94] , n_971);
  not g17524 (n_8843, n9321);
  and g17525 (\grant[94] , n_8843, n9322);
  not g17526 (n_8844, n639);
  and g17527 (n9324, n_8844, n1311);
  not g17528 (n_8845, n9324);
  and g17529 (n9325, n1316, n_8845);
  not g17530 (n_8846, n9325);
  and g17531 (n9326, n1320, n_8846);
  not g17532 (n_8847, n9326);
  and g17533 (n9327, n1324, n_8847);
  not g17534 (n_8848, n9327);
  and g17535 (n9328, n1328, n_8848);
  not g17536 (n_8849, n9328);
  and g17537 (n9329, n1332, n_8849);
  not g17538 (n_8850, n9329);
  and g17539 (n9330, n1336, n_8850);
  not g17540 (n_8851, n9330);
  and g17541 (n9331, n1340, n_8851);
  not g17542 (n_8852, n9331);
  and g17543 (n9332, n1344, n_8852);
  not g17544 (n_8853, n9332);
  and g17545 (n9333, n1348, n_8853);
  not g17546 (n_8854, n9333);
  and g17547 (n9334, n1352, n_8854);
  not g17548 (n_8855, n9334);
  and g17549 (n9335, n1356, n_8855);
  not g17550 (n_8856, n9335);
  and g17551 (n9336, n1360, n_8856);
  not g17552 (n_8857, n9336);
  and g17553 (n9337, n1364, n_8857);
  not g17554 (n_8858, n9337);
  and g17555 (n9338, n1368, n_8858);
  not g17556 (n_8859, n9338);
  and g17557 (n9339, n1372, n_8859);
  not g17558 (n_8860, n9339);
  and g17559 (n9340, n1376, n_8860);
  not g17560 (n_8861, n9340);
  and g17561 (n9341, n1380, n_8861);
  not g17562 (n_8862, n9341);
  and g17563 (n9342, n1384, n_8862);
  not g17564 (n_8863, n9342);
  and g17565 (n9343, n1388, n_8863);
  not g17566 (n_8864, n9343);
  and g17567 (n9344, n1392, n_8864);
  not g17568 (n_8865, n9344);
  and g17569 (n9345, n1396, n_8865);
  not g17570 (n_8866, n9345);
  and g17571 (n9346, n1663, n_8866);
  not g17572 (n_8867, n9346);
  and g17573 (n9347, n392, n_8867);
  not g17574 (n_8868, n9347);
  and g17575 (n9348, n396, n_8868);
  not g17576 (n_8869, n9348);
  and g17577 (n9349, n400, n_8869);
  not g17578 (n_8870, n9349);
  and g17579 (n9350, n404, n_8870);
  not g17580 (n_8871, n9350);
  and g17581 (n9351, n408, n_8871);
  not g17582 (n_8872, n9351);
  and g17583 (n9352, n412, n_8872);
  not g17584 (n_8873, n9352);
  and g17585 (n9353, n416, n_8873);
  not g17586 (n_8874, n9353);
  and g17587 (n9354, n420, n_8874);
  not g17588 (n_8875, n9354);
  and g17589 (n9355, n424, n_8875);
  not g17590 (n_8876, n9355);
  and g17591 (n9356, n428, n_8876);
  not g17592 (n_8877, n9356);
  and g17593 (n9357, n432, n_8877);
  not g17594 (n_8878, n9357);
  and g17595 (n9358, n436, n_8878);
  not g17596 (n_8879, n9358);
  and g17597 (n9359, n440, n_8879);
  not g17598 (n_8880, n9359);
  and g17599 (n9360, n444, n_8880);
  not g17600 (n_8881, n9360);
  and g17601 (n9361, n448, n_8881);
  not g17602 (n_8882, n9361);
  and g17603 (n9362, n452, n_8882);
  not g17604 (n_8883, n9362);
  and g17605 (n9363, n456, n_8883);
  not g17606 (n_8884, n9363);
  and g17607 (n9364, n460, n_8884);
  not g17608 (n_8885, n9364);
  and g17609 (n9365, n464, n_8885);
  not g17610 (n_8886, n9365);
  and g17611 (n9366, n468, n_8886);
  not g17612 (n_8887, n9366);
  and g17613 (n9367, n472, n_8887);
  not g17614 (n_8888, n9367);
  and g17615 (n9368, n476, n_8888);
  not g17616 (n_8889, n9368);
  and g17617 (n9369, n480, n_8889);
  not g17618 (n_8890, n9369);
  and g17619 (n9370, n484, n_8890);
  not g17620 (n_8891, n9370);
  and g17621 (n9371, n488, n_8891);
  not g17622 (n_8892, n9371);
  and g17623 (n9372, n492, n_8892);
  not g17624 (n_8893, n9372);
  and g17625 (n9373, n496, n_8893);
  not g17626 (n_8894, n9373);
  and g17627 (n9374, n500, n_8894);
  not g17628 (n_8895, n9374);
  and g17629 (n9375, n504, n_8895);
  not g17630 (n_8896, n9375);
  and g17631 (n9376, n508, n_8896);
  not g17632 (n_8897, n9376);
  and g17633 (n9377, n512, n_8897);
  not g17634 (n_8898, n9377);
  and g17635 (n9378, n516, n_8898);
  not g17636 (n_8899, n9378);
  and g17637 (n9379, n520, n_8899);
  not g17638 (n_8900, n9379);
  and g17639 (n9380, n524, n_8900);
  not g17640 (n_8901, n9380);
  and g17641 (n9381, n528, n_8901);
  not g17642 (n_8902, n9381);
  and g17643 (n9382, n532, n_8902);
  not g17644 (n_8903, n9382);
  and g17645 (n9383, n536, n_8903);
  not g17646 (n_8904, n9383);
  and g17647 (n9384, n540, n_8904);
  not g17648 (n_8905, n9384);
  and g17649 (n9385, n544, n_8905);
  not g17650 (n_8906, n9385);
  and g17651 (n9386, n548, n_8906);
  not g17652 (n_8907, n9386);
  and g17653 (n9387, n552, n_8907);
  not g17654 (n_8908, n9387);
  and g17655 (n9388, n556, n_8908);
  not g17656 (n_8909, n9388);
  and g17657 (n9389, n560, n_8909);
  not g17658 (n_8910, n9389);
  and g17659 (n9390, n564, n_8910);
  not g17660 (n_8911, n9390);
  and g17661 (n9391, n568, n_8911);
  not g17662 (n_8912, n9391);
  and g17663 (n9392, n572, n_8912);
  not g17664 (n_8913, n9392);
  and g17665 (n9393, n576, n_8913);
  not g17666 (n_8914, n9393);
  and g17667 (n9394, n580, n_8914);
  not g17668 (n_8915, n9394);
  and g17669 (n9395, n584, n_8915);
  not g17670 (n_8916, n9395);
  and g17671 (n9396, n588, n_8916);
  not g17672 (n_8917, n9396);
  and g17673 (n9397, n592, n_8917);
  not g17674 (n_8918, n9397);
  and g17675 (n9398, n596, n_8918);
  not g17676 (n_8919, n9398);
  and g17677 (n9399, n600, n_8919);
  not g17678 (n_8920, n9399);
  and g17679 (n9400, n604, n_8920);
  not g17680 (n_8921, n9400);
  and g17681 (n9401, n608, n_8921);
  not g17682 (n_8922, n9401);
  and g17683 (n9402, n612, n_8922);
  not g17684 (n_8923, n9402);
  and g17685 (n9403, n616, n_8923);
  not g17686 (n_8924, n9403);
  and g17687 (n9404, n620, n_8924);
  not g17688 (n_8925, n9404);
  and g17689 (n9405, n624, n_8925);
  not g17690 (n_8926, n9405);
  and g17691 (n9406, n628, n_8926);
  not g17692 (n_8927, n9406);
  and g17693 (n9407, n632, n_8927);
  and g17694 (n9408, \req[95] , n_444);
  not g17695 (n_8928, n9407);
  and g17696 (\grant[95] , n_8928, n9408);
  not g17697 (n_8929, n978);
  and g17698 (n9410, n643, n_8929);
  not g17699 (n_8930, n9410);
  and g17700 (n9411, n648, n_8930);
  not g17701 (n_8931, n9411);
  and g17702 (n9412, n652, n_8931);
  not g17703 (n_8932, n9412);
  and g17704 (n9413, n656, n_8932);
  not g17705 (n_8933, n9413);
  and g17706 (n9414, n660, n_8933);
  not g17707 (n_8934, n9414);
  and g17708 (n9415, n664, n_8934);
  not g17709 (n_8935, n9415);
  and g17710 (n9416, n668, n_8935);
  not g17711 (n_8936, n9416);
  and g17712 (n9417, n672, n_8936);
  not g17713 (n_8937, n9417);
  and g17714 (n9418, n676, n_8937);
  not g17715 (n_8938, n9418);
  and g17716 (n9419, n680, n_8938);
  not g17717 (n_8939, n9419);
  and g17718 (n9420, n684, n_8939);
  not g17719 (n_8940, n9420);
  and g17720 (n9421, n688, n_8940);
  not g17721 (n_8941, n9421);
  and g17722 (n9422, n692, n_8941);
  not g17723 (n_8942, n9422);
  and g17724 (n9423, n696, n_8942);
  not g17725 (n_8943, n9423);
  and g17726 (n9424, n700, n_8943);
  not g17727 (n_8944, n9424);
  and g17728 (n9425, n704, n_8944);
  not g17729 (n_8945, n9425);
  and g17730 (n9426, n708, n_8945);
  not g17731 (n_8946, n9426);
  and g17732 (n9427, n712, n_8946);
  not g17733 (n_8947, n9427);
  and g17734 (n9428, n716, n_8947);
  not g17735 (n_8948, n9428);
  and g17736 (n9429, n720, n_8948);
  not g17737 (n_8949, n9429);
  and g17738 (n9430, n1484, n_8949);
  not g17739 (n_8950, n9430);
  and g17740 (n9431, n1486, n_8950);
  not g17741 (n_8951, n9431);
  and g17742 (n9432, n1750, n_8951);
  not g17743 (n_8952, n9432);
  and g17744 (n9433, n731, n_8952);
  not g17745 (n_8953, n9433);
  and g17746 (n9434, n735, n_8953);
  not g17747 (n_8954, n9434);
  and g17748 (n9435, n739, n_8954);
  not g17749 (n_8955, n9435);
  and g17750 (n9436, n743, n_8955);
  not g17751 (n_8956, n9436);
  and g17752 (n9437, n747, n_8956);
  not g17753 (n_8957, n9437);
  and g17754 (n9438, n751, n_8957);
  not g17755 (n_8958, n9438);
  and g17756 (n9439, n755, n_8958);
  not g17757 (n_8959, n9439);
  and g17758 (n9440, n759, n_8959);
  not g17759 (n_8960, n9440);
  and g17760 (n9441, n763, n_8960);
  not g17761 (n_8961, n9441);
  and g17762 (n9442, n767, n_8961);
  not g17763 (n_8962, n9442);
  and g17764 (n9443, n771, n_8962);
  not g17765 (n_8963, n9443);
  and g17766 (n9444, n775, n_8963);
  not g17767 (n_8964, n9444);
  and g17768 (n9445, n779, n_8964);
  not g17769 (n_8965, n9445);
  and g17770 (n9446, n783, n_8965);
  not g17771 (n_8966, n9446);
  and g17772 (n9447, n787, n_8966);
  not g17773 (n_8967, n9447);
  and g17774 (n9448, n791, n_8967);
  not g17775 (n_8968, n9448);
  and g17776 (n9449, n795, n_8968);
  not g17777 (n_8969, n9449);
  and g17778 (n9450, n799, n_8969);
  not g17779 (n_8970, n9450);
  and g17780 (n9451, n803, n_8970);
  not g17781 (n_8971, n9451);
  and g17782 (n9452, n807, n_8971);
  not g17783 (n_8972, n9452);
  and g17784 (n9453, n811, n_8972);
  not g17785 (n_8973, n9453);
  and g17786 (n9454, n815, n_8973);
  not g17787 (n_8974, n9454);
  and g17788 (n9455, n819, n_8974);
  not g17789 (n_8975, n9455);
  and g17790 (n9456, n823, n_8975);
  not g17791 (n_8976, n9456);
  and g17792 (n9457, n827, n_8976);
  not g17793 (n_8977, n9457);
  and g17794 (n9458, n831, n_8977);
  not g17795 (n_8978, n9458);
  and g17796 (n9459, n835, n_8978);
  not g17797 (n_8979, n9459);
  and g17798 (n9460, n839, n_8979);
  not g17799 (n_8980, n9460);
  and g17800 (n9461, n843, n_8980);
  not g17801 (n_8981, n9461);
  and g17802 (n9462, n847, n_8981);
  not g17803 (n_8982, n9462);
  and g17804 (n9463, n851, n_8982);
  not g17805 (n_8983, n9463);
  and g17806 (n9464, n855, n_8983);
  not g17807 (n_8984, n9464);
  and g17808 (n9465, n859, n_8984);
  not g17809 (n_8985, n9465);
  and g17810 (n9466, n863, n_8985);
  not g17811 (n_8986, n9466);
  and g17812 (n9467, n867, n_8986);
  not g17813 (n_8987, n9467);
  and g17814 (n9468, n871, n_8987);
  not g17815 (n_8988, n9468);
  and g17816 (n9469, n875, n_8988);
  not g17817 (n_8989, n9469);
  and g17818 (n9470, n879, n_8989);
  not g17819 (n_8990, n9470);
  and g17820 (n9471, n883, n_8990);
  not g17821 (n_8991, n9471);
  and g17822 (n9472, n887, n_8991);
  not g17823 (n_8992, n9472);
  and g17824 (n9473, n891, n_8992);
  not g17825 (n_8993, n9473);
  and g17826 (n9474, n895, n_8993);
  not g17827 (n_8994, n9474);
  and g17828 (n9475, n899, n_8994);
  not g17829 (n_8995, n9475);
  and g17830 (n9476, n903, n_8995);
  not g17831 (n_8996, n9476);
  and g17832 (n9477, n907, n_8996);
  not g17833 (n_8997, n9477);
  and g17834 (n9478, n911, n_8997);
  not g17835 (n_8998, n9478);
  and g17836 (n9479, n915, n_8998);
  not g17837 (n_8999, n9479);
  and g17838 (n9480, n919, n_8999);
  not g17839 (n_9000, n9480);
  and g17840 (n9481, n923, n_9000);
  not g17841 (n_9001, n9481);
  and g17842 (n9482, n927, n_9001);
  not g17843 (n_9002, n9482);
  and g17844 (n9483, n931, n_9002);
  not g17845 (n_9003, n9483);
  and g17846 (n9484, n935, n_9003);
  not g17847 (n_9004, n9484);
  and g17848 (n9485, n939, n_9004);
  not g17849 (n_9005, n9485);
  and g17850 (n9486, n943, n_9005);
  not g17851 (n_9006, n9486);
  and g17852 (n9487, n947, n_9006);
  not g17853 (n_9007, n9487);
  and g17854 (n9488, n951, n_9007);
  not g17855 (n_9008, n9488);
  and g17856 (n9489, n955, n_9008);
  not g17857 (n_9009, n9489);
  and g17858 (n9490, n959, n_9009);
  not g17859 (n_9010, n9490);
  and g17860 (n9491, n963, n_9010);
  not g17861 (n_9011, n9491);
  and g17862 (n9492, n967, n_9011);
  not g17863 (n_9012, n9492);
  and g17864 (n9493, n971, n_9012);
  and g17865 (n9494, \req[96] , n_785);
  not g17866 (n_9013, n9493);
  and g17867 (\grant[96] , n_9013, n9494);
  not g17868 (n_9014, n1315);
  and g17869 (n9496, n982, n_9014);
  not g17870 (n_9015, n9496);
  and g17871 (n9497, n987, n_9015);
  not g17872 (n_9016, n9497);
  and g17873 (n9498, n991, n_9016);
  not g17874 (n_9017, n9498);
  and g17875 (n9499, n995, n_9017);
  not g17876 (n_9018, n9499);
  and g17877 (n9500, n999, n_9018);
  not g17878 (n_9019, n9500);
  and g17879 (n9501, n1003, n_9019);
  not g17880 (n_9020, n9501);
  and g17881 (n9502, n1007, n_9020);
  not g17882 (n_9021, n9502);
  and g17883 (n9503, n1011, n_9021);
  not g17884 (n_9022, n9503);
  and g17885 (n9504, n1015, n_9022);
  not g17886 (n_9023, n9504);
  and g17887 (n9505, n1019, n_9023);
  not g17888 (n_9024, n9505);
  and g17889 (n9506, n1023, n_9024);
  not g17890 (n_9025, n9506);
  and g17891 (n9507, n1027, n_9025);
  not g17892 (n_9026, n9507);
  and g17893 (n9508, n1031, n_9026);
  not g17894 (n_9027, n9508);
  and g17895 (n9509, n1035, n_9027);
  not g17896 (n_9028, n9509);
  and g17897 (n9510, n1039, n_9028);
  not g17898 (n_9029, n9510);
  and g17899 (n9511, n1043, n_9029);
  not g17900 (n_9030, n9511);
  and g17901 (n9512, n1047, n_9030);
  not g17902 (n_9031, n9512);
  and g17903 (n9513, n1051, n_9031);
  not g17904 (n_9032, n9513);
  and g17905 (n9514, n1055, n_9032);
  not g17906 (n_9033, n9514);
  and g17907 (n9515, n1059, n_9033);
  not g17908 (n_9034, n9515);
  and g17909 (n9516, n1574, n_9034);
  not g17910 (n_9035, n9516);
  and g17911 (n9517, n1576, n_9035);
  not g17912 (n_9036, n9517);
  and g17913 (n9518, n1837, n_9036);
  not g17914 (n_9037, n9518);
  and g17915 (n9519, n1068, n_9037);
  not g17916 (n_9038, n9519);
  and g17917 (n9520, n1072, n_9038);
  not g17918 (n_9039, n9520);
  and g17919 (n9521, n1076, n_9039);
  not g17920 (n_9040, n9521);
  and g17921 (n9522, n1080, n_9040);
  not g17922 (n_9041, n9522);
  and g17923 (n9523, n1084, n_9041);
  not g17924 (n_9042, n9523);
  and g17925 (n9524, n1088, n_9042);
  not g17926 (n_9043, n9524);
  and g17927 (n9525, n1092, n_9043);
  not g17928 (n_9044, n9525);
  and g17929 (n9526, n1096, n_9044);
  not g17930 (n_9045, n9526);
  and g17931 (n9527, n1100, n_9045);
  not g17932 (n_9046, n9527);
  and g17933 (n9528, n1104, n_9046);
  not g17934 (n_9047, n9528);
  and g17935 (n9529, n1108, n_9047);
  not g17936 (n_9048, n9529);
  and g17937 (n9530, n1112, n_9048);
  not g17938 (n_9049, n9530);
  and g17939 (n9531, n1116, n_9049);
  not g17940 (n_9050, n9531);
  and g17941 (n9532, n1120, n_9050);
  not g17942 (n_9051, n9532);
  and g17943 (n9533, n1124, n_9051);
  not g17944 (n_9052, n9533);
  and g17945 (n9534, n1128, n_9052);
  not g17946 (n_9053, n9534);
  and g17947 (n9535, n1132, n_9053);
  not g17948 (n_9054, n9535);
  and g17949 (n9536, n1136, n_9054);
  not g17950 (n_9055, n9536);
  and g17951 (n9537, n1140, n_9055);
  not g17952 (n_9056, n9537);
  and g17953 (n9538, n1144, n_9056);
  not g17954 (n_9057, n9538);
  and g17955 (n9539, n1148, n_9057);
  not g17956 (n_9058, n9539);
  and g17957 (n9540, n1152, n_9058);
  not g17958 (n_9059, n9540);
  and g17959 (n9541, n1156, n_9059);
  not g17960 (n_9060, n9541);
  and g17961 (n9542, n1160, n_9060);
  not g17962 (n_9061, n9542);
  and g17963 (n9543, n1164, n_9061);
  not g17964 (n_9062, n9543);
  and g17965 (n9544, n1168, n_9062);
  not g17966 (n_9063, n9544);
  and g17967 (n9545, n1172, n_9063);
  not g17968 (n_9064, n9545);
  and g17969 (n9546, n1176, n_9064);
  not g17970 (n_9065, n9546);
  and g17971 (n9547, n1180, n_9065);
  not g17972 (n_9066, n9547);
  and g17973 (n9548, n1184, n_9066);
  not g17974 (n_9067, n9548);
  and g17975 (n9549, n1188, n_9067);
  not g17976 (n_9068, n9549);
  and g17977 (n9550, n1192, n_9068);
  not g17978 (n_9069, n9550);
  and g17979 (n9551, n1196, n_9069);
  not g17980 (n_9070, n9551);
  and g17981 (n9552, n1200, n_9070);
  not g17982 (n_9071, n9552);
  and g17983 (n9553, n1204, n_9071);
  not g17984 (n_9072, n9553);
  and g17985 (n9554, n1208, n_9072);
  not g17986 (n_9073, n9554);
  and g17987 (n9555, n1212, n_9073);
  not g17988 (n_9074, n9555);
  and g17989 (n9556, n1216, n_9074);
  not g17990 (n_9075, n9556);
  and g17991 (n9557, n1220, n_9075);
  not g17992 (n_9076, n9557);
  and g17993 (n9558, n1224, n_9076);
  not g17994 (n_9077, n9558);
  and g17995 (n9559, n1228, n_9077);
  not g17996 (n_9078, n9559);
  and g17997 (n9560, n1232, n_9078);
  not g17998 (n_9079, n9560);
  and g17999 (n9561, n1236, n_9079);
  not g18000 (n_9080, n9561);
  and g18001 (n9562, n1240, n_9080);
  not g18002 (n_9081, n9562);
  and g18003 (n9563, n1244, n_9081);
  not g18004 (n_9082, n9563);
  and g18005 (n9564, n1248, n_9082);
  not g18006 (n_9083, n9564);
  and g18007 (n9565, n1252, n_9083);
  not g18008 (n_9084, n9565);
  and g18009 (n9566, n1256, n_9084);
  not g18010 (n_9085, n9566);
  and g18011 (n9567, n1260, n_9085);
  not g18012 (n_9086, n9567);
  and g18013 (n9568, n1264, n_9086);
  not g18014 (n_9087, n9568);
  and g18015 (n9569, n1268, n_9087);
  not g18016 (n_9088, n9569);
  and g18017 (n9570, n1272, n_9088);
  not g18018 (n_9089, n9570);
  and g18019 (n9571, n1276, n_9089);
  not g18020 (n_9090, n9571);
  and g18021 (n9572, n1280, n_9090);
  not g18022 (n_9091, n9572);
  and g18023 (n9573, n1284, n_9091);
  not g18024 (n_9092, n9573);
  and g18025 (n9574, n1288, n_9092);
  not g18026 (n_9093, n9574);
  and g18027 (n9575, n1292, n_9093);
  not g18028 (n_9094, n9575);
  and g18029 (n9576, n1296, n_9094);
  not g18030 (n_9095, n9576);
  and g18031 (n9577, n1300, n_9095);
  not g18032 (n_9096, n9577);
  and g18033 (n9578, n1304, n_9096);
  not g18034 (n_9097, n9578);
  and g18035 (n9579, n1308, n_9097);
  and g18036 (n9580, \req[97] , n_975);
  not g18037 (n_9098, n9579);
  and g18038 (\grant[97] , n_9098, n9580);
  not g18039 (n_9099, n647);
  and g18040 (n9582, n_9099, n1319);
  not g18041 (n_9100, n9582);
  and g18042 (n9583, n1324, n_9100);
  not g18043 (n_9101, n9583);
  and g18044 (n9584, n1328, n_9101);
  not g18045 (n_9102, n9584);
  and g18046 (n9585, n1332, n_9102);
  not g18047 (n_9103, n9585);
  and g18048 (n9586, n1336, n_9103);
  not g18049 (n_9104, n9586);
  and g18050 (n9587, n1340, n_9104);
  not g18051 (n_9105, n9587);
  and g18052 (n9588, n1344, n_9105);
  not g18053 (n_9106, n9588);
  and g18054 (n9589, n1348, n_9106);
  not g18055 (n_9107, n9589);
  and g18056 (n9590, n1352, n_9107);
  not g18057 (n_9108, n9590);
  and g18058 (n9591, n1356, n_9108);
  not g18059 (n_9109, n9591);
  and g18060 (n9592, n1360, n_9109);
  not g18061 (n_9110, n9592);
  and g18062 (n9593, n1364, n_9110);
  not g18063 (n_9111, n9593);
  and g18064 (n9594, n1368, n_9111);
  not g18065 (n_9112, n9594);
  and g18066 (n9595, n1372, n_9112);
  not g18067 (n_9113, n9595);
  and g18068 (n9596, n1376, n_9113);
  not g18069 (n_9114, n9596);
  and g18070 (n9597, n1380, n_9114);
  not g18071 (n_9115, n9597);
  and g18072 (n9598, n1384, n_9115);
  not g18073 (n_9116, n9598);
  and g18074 (n9599, n1388, n_9116);
  not g18075 (n_9117, n9599);
  and g18076 (n9600, n1392, n_9117);
  not g18077 (n_9118, n9600);
  and g18078 (n9601, n1396, n_9118);
  not g18079 (n_9119, n9601);
  and g18080 (n9602, n1663, n_9119);
  not g18081 (n_9120, n9602);
  and g18082 (n9603, n392, n_9120);
  not g18083 (n_9121, n9603);
  and g18084 (n9604, n396, n_9121);
  not g18085 (n_9122, n9604);
  and g18086 (n9605, n400, n_9122);
  not g18087 (n_9123, n9605);
  and g18088 (n9606, n404, n_9123);
  not g18089 (n_9124, n9606);
  and g18090 (n9607, n408, n_9124);
  not g18091 (n_9125, n9607);
  and g18092 (n9608, n412, n_9125);
  not g18093 (n_9126, n9608);
  and g18094 (n9609, n416, n_9126);
  not g18095 (n_9127, n9609);
  and g18096 (n9610, n420, n_9127);
  not g18097 (n_9128, n9610);
  and g18098 (n9611, n424, n_9128);
  not g18099 (n_9129, n9611);
  and g18100 (n9612, n428, n_9129);
  not g18101 (n_9130, n9612);
  and g18102 (n9613, n432, n_9130);
  not g18103 (n_9131, n9613);
  and g18104 (n9614, n436, n_9131);
  not g18105 (n_9132, n9614);
  and g18106 (n9615, n440, n_9132);
  not g18107 (n_9133, n9615);
  and g18108 (n9616, n444, n_9133);
  not g18109 (n_9134, n9616);
  and g18110 (n9617, n448, n_9134);
  not g18111 (n_9135, n9617);
  and g18112 (n9618, n452, n_9135);
  not g18113 (n_9136, n9618);
  and g18114 (n9619, n456, n_9136);
  not g18115 (n_9137, n9619);
  and g18116 (n9620, n460, n_9137);
  not g18117 (n_9138, n9620);
  and g18118 (n9621, n464, n_9138);
  not g18119 (n_9139, n9621);
  and g18120 (n9622, n468, n_9139);
  not g18121 (n_9140, n9622);
  and g18122 (n9623, n472, n_9140);
  not g18123 (n_9141, n9623);
  and g18124 (n9624, n476, n_9141);
  not g18125 (n_9142, n9624);
  and g18126 (n9625, n480, n_9142);
  not g18127 (n_9143, n9625);
  and g18128 (n9626, n484, n_9143);
  not g18129 (n_9144, n9626);
  and g18130 (n9627, n488, n_9144);
  not g18131 (n_9145, n9627);
  and g18132 (n9628, n492, n_9145);
  not g18133 (n_9146, n9628);
  and g18134 (n9629, n496, n_9146);
  not g18135 (n_9147, n9629);
  and g18136 (n9630, n500, n_9147);
  not g18137 (n_9148, n9630);
  and g18138 (n9631, n504, n_9148);
  not g18139 (n_9149, n9631);
  and g18140 (n9632, n508, n_9149);
  not g18141 (n_9150, n9632);
  and g18142 (n9633, n512, n_9150);
  not g18143 (n_9151, n9633);
  and g18144 (n9634, n516, n_9151);
  not g18145 (n_9152, n9634);
  and g18146 (n9635, n520, n_9152);
  not g18147 (n_9153, n9635);
  and g18148 (n9636, n524, n_9153);
  not g18149 (n_9154, n9636);
  and g18150 (n9637, n528, n_9154);
  not g18151 (n_9155, n9637);
  and g18152 (n9638, n532, n_9155);
  not g18153 (n_9156, n9638);
  and g18154 (n9639, n536, n_9156);
  not g18155 (n_9157, n9639);
  and g18156 (n9640, n540, n_9157);
  not g18157 (n_9158, n9640);
  and g18158 (n9641, n544, n_9158);
  not g18159 (n_9159, n9641);
  and g18160 (n9642, n548, n_9159);
  not g18161 (n_9160, n9642);
  and g18162 (n9643, n552, n_9160);
  not g18163 (n_9161, n9643);
  and g18164 (n9644, n556, n_9161);
  not g18165 (n_9162, n9644);
  and g18166 (n9645, n560, n_9162);
  not g18167 (n_9163, n9645);
  and g18168 (n9646, n564, n_9163);
  not g18169 (n_9164, n9646);
  and g18170 (n9647, n568, n_9164);
  not g18171 (n_9165, n9647);
  and g18172 (n9648, n572, n_9165);
  not g18173 (n_9166, n9648);
  and g18174 (n9649, n576, n_9166);
  not g18175 (n_9167, n9649);
  and g18176 (n9650, n580, n_9167);
  not g18177 (n_9168, n9650);
  and g18178 (n9651, n584, n_9168);
  not g18179 (n_9169, n9651);
  and g18180 (n9652, n588, n_9169);
  not g18181 (n_9170, n9652);
  and g18182 (n9653, n592, n_9170);
  not g18183 (n_9171, n9653);
  and g18184 (n9654, n596, n_9171);
  not g18185 (n_9172, n9654);
  and g18186 (n9655, n600, n_9172);
  not g18187 (n_9173, n9655);
  and g18188 (n9656, n604, n_9173);
  not g18189 (n_9174, n9656);
  and g18190 (n9657, n608, n_9174);
  not g18191 (n_9175, n9657);
  and g18192 (n9658, n612, n_9175);
  not g18193 (n_9176, n9658);
  and g18194 (n9659, n616, n_9176);
  not g18195 (n_9177, n9659);
  and g18196 (n9660, n620, n_9177);
  not g18197 (n_9178, n9660);
  and g18198 (n9661, n624, n_9178);
  not g18199 (n_9179, n9661);
  and g18200 (n9662, n628, n_9179);
  not g18201 (n_9180, n9662);
  and g18202 (n9663, n632, n_9180);
  not g18203 (n_9181, n9663);
  and g18204 (n9664, n636, n_9181);
  not g18205 (n_9182, n9664);
  and g18206 (n9665, n640, n_9182);
  and g18207 (n9666, \req[98] , n_458);
  not g18208 (n_9183, n9665);
  and g18209 (\grant[98] , n_9183, n9666);
  not g18210 (n_9184, n986);
  and g18211 (n9668, n651, n_9184);
  not g18212 (n_9185, n9668);
  and g18213 (n9669, n656, n_9185);
  not g18214 (n_9186, n9669);
  and g18215 (n9670, n660, n_9186);
  not g18216 (n_9187, n9670);
  and g18217 (n9671, n664, n_9187);
  not g18218 (n_9188, n9671);
  and g18219 (n9672, n668, n_9188);
  not g18220 (n_9189, n9672);
  and g18221 (n9673, n672, n_9189);
  not g18222 (n_9190, n9673);
  and g18223 (n9674, n676, n_9190);
  not g18224 (n_9191, n9674);
  and g18225 (n9675, n680, n_9191);
  not g18226 (n_9192, n9675);
  and g18227 (n9676, n684, n_9192);
  not g18228 (n_9193, n9676);
  and g18229 (n9677, n688, n_9193);
  not g18230 (n_9194, n9677);
  and g18231 (n9678, n692, n_9194);
  not g18232 (n_9195, n9678);
  and g18233 (n9679, n696, n_9195);
  not g18234 (n_9196, n9679);
  and g18235 (n9680, n700, n_9196);
  not g18236 (n_9197, n9680);
  and g18237 (n9681, n704, n_9197);
  not g18238 (n_9198, n9681);
  and g18239 (n9682, n708, n_9198);
  not g18240 (n_9199, n9682);
  and g18241 (n9683, n712, n_9199);
  not g18242 (n_9200, n9683);
  and g18243 (n9684, n716, n_9200);
  not g18244 (n_9201, n9684);
  and g18245 (n9685, n720, n_9201);
  not g18246 (n_9202, n9685);
  and g18247 (n9686, n1484, n_9202);
  not g18248 (n_9203, n9686);
  and g18249 (n9687, n1486, n_9203);
  not g18250 (n_9204, n9687);
  and g18251 (n9688, n1750, n_9204);
  not g18252 (n_9205, n9688);
  and g18253 (n9689, n731, n_9205);
  not g18254 (n_9206, n9689);
  and g18255 (n9690, n735, n_9206);
  not g18256 (n_9207, n9690);
  and g18257 (n9691, n739, n_9207);
  not g18258 (n_9208, n9691);
  and g18259 (n9692, n743, n_9208);
  not g18260 (n_9209, n9692);
  and g18261 (n9693, n747, n_9209);
  not g18262 (n_9210, n9693);
  and g18263 (n9694, n751, n_9210);
  not g18264 (n_9211, n9694);
  and g18265 (n9695, n755, n_9211);
  not g18266 (n_9212, n9695);
  and g18267 (n9696, n759, n_9212);
  not g18268 (n_9213, n9696);
  and g18269 (n9697, n763, n_9213);
  not g18270 (n_9214, n9697);
  and g18271 (n9698, n767, n_9214);
  not g18272 (n_9215, n9698);
  and g18273 (n9699, n771, n_9215);
  not g18274 (n_9216, n9699);
  and g18275 (n9700, n775, n_9216);
  not g18276 (n_9217, n9700);
  and g18277 (n9701, n779, n_9217);
  not g18278 (n_9218, n9701);
  and g18279 (n9702, n783, n_9218);
  not g18280 (n_9219, n9702);
  and g18281 (n9703, n787, n_9219);
  not g18282 (n_9220, n9703);
  and g18283 (n9704, n791, n_9220);
  not g18284 (n_9221, n9704);
  and g18285 (n9705, n795, n_9221);
  not g18286 (n_9222, n9705);
  and g18287 (n9706, n799, n_9222);
  not g18288 (n_9223, n9706);
  and g18289 (n9707, n803, n_9223);
  not g18290 (n_9224, n9707);
  and g18291 (n9708, n807, n_9224);
  not g18292 (n_9225, n9708);
  and g18293 (n9709, n811, n_9225);
  not g18294 (n_9226, n9709);
  and g18295 (n9710, n815, n_9226);
  not g18296 (n_9227, n9710);
  and g18297 (n9711, n819, n_9227);
  not g18298 (n_9228, n9711);
  and g18299 (n9712, n823, n_9228);
  not g18300 (n_9229, n9712);
  and g18301 (n9713, n827, n_9229);
  not g18302 (n_9230, n9713);
  and g18303 (n9714, n831, n_9230);
  not g18304 (n_9231, n9714);
  and g18305 (n9715, n835, n_9231);
  not g18306 (n_9232, n9715);
  and g18307 (n9716, n839, n_9232);
  not g18308 (n_9233, n9716);
  and g18309 (n9717, n843, n_9233);
  not g18310 (n_9234, n9717);
  and g18311 (n9718, n847, n_9234);
  not g18312 (n_9235, n9718);
  and g18313 (n9719, n851, n_9235);
  not g18314 (n_9236, n9719);
  and g18315 (n9720, n855, n_9236);
  not g18316 (n_9237, n9720);
  and g18317 (n9721, n859, n_9237);
  not g18318 (n_9238, n9721);
  and g18319 (n9722, n863, n_9238);
  not g18320 (n_9239, n9722);
  and g18321 (n9723, n867, n_9239);
  not g18322 (n_9240, n9723);
  and g18323 (n9724, n871, n_9240);
  not g18324 (n_9241, n9724);
  and g18325 (n9725, n875, n_9241);
  not g18326 (n_9242, n9725);
  and g18327 (n9726, n879, n_9242);
  not g18328 (n_9243, n9726);
  and g18329 (n9727, n883, n_9243);
  not g18330 (n_9244, n9727);
  and g18331 (n9728, n887, n_9244);
  not g18332 (n_9245, n9728);
  and g18333 (n9729, n891, n_9245);
  not g18334 (n_9246, n9729);
  and g18335 (n9730, n895, n_9246);
  not g18336 (n_9247, n9730);
  and g18337 (n9731, n899, n_9247);
  not g18338 (n_9248, n9731);
  and g18339 (n9732, n903, n_9248);
  not g18340 (n_9249, n9732);
  and g18341 (n9733, n907, n_9249);
  not g18342 (n_9250, n9733);
  and g18343 (n9734, n911, n_9250);
  not g18344 (n_9251, n9734);
  and g18345 (n9735, n915, n_9251);
  not g18346 (n_9252, n9735);
  and g18347 (n9736, n919, n_9252);
  not g18348 (n_9253, n9736);
  and g18349 (n9737, n923, n_9253);
  not g18350 (n_9254, n9737);
  and g18351 (n9738, n927, n_9254);
  not g18352 (n_9255, n9738);
  and g18353 (n9739, n931, n_9255);
  not g18354 (n_9256, n9739);
  and g18355 (n9740, n935, n_9256);
  not g18356 (n_9257, n9740);
  and g18357 (n9741, n939, n_9257);
  not g18358 (n_9258, n9741);
  and g18359 (n9742, n943, n_9258);
  not g18360 (n_9259, n9742);
  and g18361 (n9743, n947, n_9259);
  not g18362 (n_9260, n9743);
  and g18363 (n9744, n951, n_9260);
  not g18364 (n_9261, n9744);
  and g18365 (n9745, n955, n_9261);
  not g18366 (n_9262, n9745);
  and g18367 (n9746, n959, n_9262);
  not g18368 (n_9263, n9746);
  and g18369 (n9747, n963, n_9263);
  not g18370 (n_9264, n9747);
  and g18371 (n9748, n967, n_9264);
  not g18372 (n_9265, n9748);
  and g18373 (n9749, n971, n_9265);
  not g18374 (n_9266, n9749);
  and g18375 (n9750, n975, n_9266);
  not g18376 (n_9267, n9750);
  and g18377 (n9751, n979, n_9267);
  and g18378 (n9752, \req[99] , n_791);
  not g18379 (n_9268, n9751);
  and g18380 (\grant[99] , n_9268, n9752);
  not g18381 (n_9269, n1323);
  and g18382 (n9754, n990, n_9269);
  not g18383 (n_9270, n9754);
  and g18384 (n9755, n995, n_9270);
  not g18385 (n_9271, n9755);
  and g18386 (n9756, n999, n_9271);
  not g18387 (n_9272, n9756);
  and g18388 (n9757, n1003, n_9272);
  not g18389 (n_9273, n9757);
  and g18390 (n9758, n1007, n_9273);
  not g18391 (n_9274, n9758);
  and g18392 (n9759, n1011, n_9274);
  not g18393 (n_9275, n9759);
  and g18394 (n9760, n1015, n_9275);
  not g18395 (n_9276, n9760);
  and g18396 (n9761, n1019, n_9276);
  not g18397 (n_9277, n9761);
  and g18398 (n9762, n1023, n_9277);
  not g18399 (n_9278, n9762);
  and g18400 (n9763, n1027, n_9278);
  not g18401 (n_9279, n9763);
  and g18402 (n9764, n1031, n_9279);
  not g18403 (n_9280, n9764);
  and g18404 (n9765, n1035, n_9280);
  not g18405 (n_9281, n9765);
  and g18406 (n9766, n1039, n_9281);
  not g18407 (n_9282, n9766);
  and g18408 (n9767, n1043, n_9282);
  not g18409 (n_9283, n9767);
  and g18410 (n9768, n1047, n_9283);
  not g18411 (n_9284, n9768);
  and g18412 (n9769, n1051, n_9284);
  not g18413 (n_9285, n9769);
  and g18414 (n9770, n1055, n_9285);
  not g18415 (n_9286, n9770);
  and g18416 (n9771, n1059, n_9286);
  not g18417 (n_9287, n9771);
  and g18418 (n9772, n1574, n_9287);
  not g18419 (n_9288, n9772);
  and g18420 (n9773, n1576, n_9288);
  not g18421 (n_9289, n9773);
  and g18422 (n9774, n1837, n_9289);
  not g18423 (n_9290, n9774);
  and g18424 (n9775, n1068, n_9290);
  not g18425 (n_9291, n9775);
  and g18426 (n9776, n1072, n_9291);
  not g18427 (n_9292, n9776);
  and g18428 (n9777, n1076, n_9292);
  not g18429 (n_9293, n9777);
  and g18430 (n9778, n1080, n_9293);
  not g18431 (n_9294, n9778);
  and g18432 (n9779, n1084, n_9294);
  not g18433 (n_9295, n9779);
  and g18434 (n9780, n1088, n_9295);
  not g18435 (n_9296, n9780);
  and g18436 (n9781, n1092, n_9296);
  not g18437 (n_9297, n9781);
  and g18438 (n9782, n1096, n_9297);
  not g18439 (n_9298, n9782);
  and g18440 (n9783, n1100, n_9298);
  not g18441 (n_9299, n9783);
  and g18442 (n9784, n1104, n_9299);
  not g18443 (n_9300, n9784);
  and g18444 (n9785, n1108, n_9300);
  not g18445 (n_9301, n9785);
  and g18446 (n9786, n1112, n_9301);
  not g18447 (n_9302, n9786);
  and g18448 (n9787, n1116, n_9302);
  not g18449 (n_9303, n9787);
  and g18450 (n9788, n1120, n_9303);
  not g18451 (n_9304, n9788);
  and g18452 (n9789, n1124, n_9304);
  not g18453 (n_9305, n9789);
  and g18454 (n9790, n1128, n_9305);
  not g18455 (n_9306, n9790);
  and g18456 (n9791, n1132, n_9306);
  not g18457 (n_9307, n9791);
  and g18458 (n9792, n1136, n_9307);
  not g18459 (n_9308, n9792);
  and g18460 (n9793, n1140, n_9308);
  not g18461 (n_9309, n9793);
  and g18462 (n9794, n1144, n_9309);
  not g18463 (n_9310, n9794);
  and g18464 (n9795, n1148, n_9310);
  not g18465 (n_9311, n9795);
  and g18466 (n9796, n1152, n_9311);
  not g18467 (n_9312, n9796);
  and g18468 (n9797, n1156, n_9312);
  not g18469 (n_9313, n9797);
  and g18470 (n9798, n1160, n_9313);
  not g18471 (n_9314, n9798);
  and g18472 (n9799, n1164, n_9314);
  not g18473 (n_9315, n9799);
  and g18474 (n9800, n1168, n_9315);
  not g18475 (n_9316, n9800);
  and g18476 (n9801, n1172, n_9316);
  not g18477 (n_9317, n9801);
  and g18478 (n9802, n1176, n_9317);
  not g18479 (n_9318, n9802);
  and g18480 (n9803, n1180, n_9318);
  not g18481 (n_9319, n9803);
  and g18482 (n9804, n1184, n_9319);
  not g18483 (n_9320, n9804);
  and g18484 (n9805, n1188, n_9320);
  not g18485 (n_9321, n9805);
  and g18486 (n9806, n1192, n_9321);
  not g18487 (n_9322, n9806);
  and g18488 (n9807, n1196, n_9322);
  not g18489 (n_9323, n9807);
  and g18490 (n9808, n1200, n_9323);
  not g18491 (n_9324, n9808);
  and g18492 (n9809, n1204, n_9324);
  not g18493 (n_9325, n9809);
  and g18494 (n9810, n1208, n_9325);
  not g18495 (n_9326, n9810);
  and g18496 (n9811, n1212, n_9326);
  not g18497 (n_9327, n9811);
  and g18498 (n9812, n1216, n_9327);
  not g18499 (n_9328, n9812);
  and g18500 (n9813, n1220, n_9328);
  not g18501 (n_9329, n9813);
  and g18502 (n9814, n1224, n_9329);
  not g18503 (n_9330, n9814);
  and g18504 (n9815, n1228, n_9330);
  not g18505 (n_9331, n9815);
  and g18506 (n9816, n1232, n_9331);
  not g18507 (n_9332, n9816);
  and g18508 (n9817, n1236, n_9332);
  not g18509 (n_9333, n9817);
  and g18510 (n9818, n1240, n_9333);
  not g18511 (n_9334, n9818);
  and g18512 (n9819, n1244, n_9334);
  not g18513 (n_9335, n9819);
  and g18514 (n9820, n1248, n_9335);
  not g18515 (n_9336, n9820);
  and g18516 (n9821, n1252, n_9336);
  not g18517 (n_9337, n9821);
  and g18518 (n9822, n1256, n_9337);
  not g18519 (n_9338, n9822);
  and g18520 (n9823, n1260, n_9338);
  not g18521 (n_9339, n9823);
  and g18522 (n9824, n1264, n_9339);
  not g18523 (n_9340, n9824);
  and g18524 (n9825, n1268, n_9340);
  not g18525 (n_9341, n9825);
  and g18526 (n9826, n1272, n_9341);
  not g18527 (n_9342, n9826);
  and g18528 (n9827, n1276, n_9342);
  not g18529 (n_9343, n9827);
  and g18530 (n9828, n1280, n_9343);
  not g18531 (n_9344, n9828);
  and g18532 (n9829, n1284, n_9344);
  not g18533 (n_9345, n9829);
  and g18534 (n9830, n1288, n_9345);
  not g18535 (n_9346, n9830);
  and g18536 (n9831, n1292, n_9346);
  not g18537 (n_9347, n9831);
  and g18538 (n9832, n1296, n_9347);
  not g18539 (n_9348, n9832);
  and g18540 (n9833, n1300, n_9348);
  not g18541 (n_9349, n9833);
  and g18542 (n9834, n1304, n_9349);
  not g18543 (n_9350, n9834);
  and g18544 (n9835, n1308, n_9350);
  not g18545 (n_9351, n9835);
  and g18546 (n9836, n1312, n_9351);
  not g18547 (n_9352, n9836);
  and g18548 (n9837, n1316, n_9352);
  and g18549 (n9838, \req[100] , n_979);
  not g18550 (n_9353, n9837);
  and g18551 (\grant[100] , n_9353, n9838);
  not g18552 (n_9354, n655);
  and g18553 (n9840, n_9354, n1327);
  not g18554 (n_9355, n9840);
  and g18555 (n9841, n1332, n_9355);
  not g18556 (n_9356, n9841);
  and g18557 (n9842, n1336, n_9356);
  not g18558 (n_9357, n9842);
  and g18559 (n9843, n1340, n_9357);
  not g18560 (n_9358, n9843);
  and g18561 (n9844, n1344, n_9358);
  not g18562 (n_9359, n9844);
  and g18563 (n9845, n1348, n_9359);
  not g18564 (n_9360, n9845);
  and g18565 (n9846, n1352, n_9360);
  not g18566 (n_9361, n9846);
  and g18567 (n9847, n1356, n_9361);
  not g18568 (n_9362, n9847);
  and g18569 (n9848, n1360, n_9362);
  not g18570 (n_9363, n9848);
  and g18571 (n9849, n1364, n_9363);
  not g18572 (n_9364, n9849);
  and g18573 (n9850, n1368, n_9364);
  not g18574 (n_9365, n9850);
  and g18575 (n9851, n1372, n_9365);
  not g18576 (n_9366, n9851);
  and g18577 (n9852, n1376, n_9366);
  not g18578 (n_9367, n9852);
  and g18579 (n9853, n1380, n_9367);
  not g18580 (n_9368, n9853);
  and g18581 (n9854, n1384, n_9368);
  not g18582 (n_9369, n9854);
  and g18583 (n9855, n1388, n_9369);
  not g18584 (n_9370, n9855);
  and g18585 (n9856, n1392, n_9370);
  not g18586 (n_9371, n9856);
  and g18587 (n9857, n1396, n_9371);
  not g18588 (n_9372, n9857);
  and g18589 (n9858, n1663, n_9372);
  not g18590 (n_9373, n9858);
  and g18591 (n9859, n392, n_9373);
  not g18592 (n_9374, n9859);
  and g18593 (n9860, n396, n_9374);
  not g18594 (n_9375, n9860);
  and g18595 (n9861, n400, n_9375);
  not g18596 (n_9376, n9861);
  and g18597 (n9862, n404, n_9376);
  not g18598 (n_9377, n9862);
  and g18599 (n9863, n408, n_9377);
  not g18600 (n_9378, n9863);
  and g18601 (n9864, n412, n_9378);
  not g18602 (n_9379, n9864);
  and g18603 (n9865, n416, n_9379);
  not g18604 (n_9380, n9865);
  and g18605 (n9866, n420, n_9380);
  not g18606 (n_9381, n9866);
  and g18607 (n9867, n424, n_9381);
  not g18608 (n_9382, n9867);
  and g18609 (n9868, n428, n_9382);
  not g18610 (n_9383, n9868);
  and g18611 (n9869, n432, n_9383);
  not g18612 (n_9384, n9869);
  and g18613 (n9870, n436, n_9384);
  not g18614 (n_9385, n9870);
  and g18615 (n9871, n440, n_9385);
  not g18616 (n_9386, n9871);
  and g18617 (n9872, n444, n_9386);
  not g18618 (n_9387, n9872);
  and g18619 (n9873, n448, n_9387);
  not g18620 (n_9388, n9873);
  and g18621 (n9874, n452, n_9388);
  not g18622 (n_9389, n9874);
  and g18623 (n9875, n456, n_9389);
  not g18624 (n_9390, n9875);
  and g18625 (n9876, n460, n_9390);
  not g18626 (n_9391, n9876);
  and g18627 (n9877, n464, n_9391);
  not g18628 (n_9392, n9877);
  and g18629 (n9878, n468, n_9392);
  not g18630 (n_9393, n9878);
  and g18631 (n9879, n472, n_9393);
  not g18632 (n_9394, n9879);
  and g18633 (n9880, n476, n_9394);
  not g18634 (n_9395, n9880);
  and g18635 (n9881, n480, n_9395);
  not g18636 (n_9396, n9881);
  and g18637 (n9882, n484, n_9396);
  not g18638 (n_9397, n9882);
  and g18639 (n9883, n488, n_9397);
  not g18640 (n_9398, n9883);
  and g18641 (n9884, n492, n_9398);
  not g18642 (n_9399, n9884);
  and g18643 (n9885, n496, n_9399);
  not g18644 (n_9400, n9885);
  and g18645 (n9886, n500, n_9400);
  not g18646 (n_9401, n9886);
  and g18647 (n9887, n504, n_9401);
  not g18648 (n_9402, n9887);
  and g18649 (n9888, n508, n_9402);
  not g18650 (n_9403, n9888);
  and g18651 (n9889, n512, n_9403);
  not g18652 (n_9404, n9889);
  and g18653 (n9890, n516, n_9404);
  not g18654 (n_9405, n9890);
  and g18655 (n9891, n520, n_9405);
  not g18656 (n_9406, n9891);
  and g18657 (n9892, n524, n_9406);
  not g18658 (n_9407, n9892);
  and g18659 (n9893, n528, n_9407);
  not g18660 (n_9408, n9893);
  and g18661 (n9894, n532, n_9408);
  not g18662 (n_9409, n9894);
  and g18663 (n9895, n536, n_9409);
  not g18664 (n_9410, n9895);
  and g18665 (n9896, n540, n_9410);
  not g18666 (n_9411, n9896);
  and g18667 (n9897, n544, n_9411);
  not g18668 (n_9412, n9897);
  and g18669 (n9898, n548, n_9412);
  not g18670 (n_9413, n9898);
  and g18671 (n9899, n552, n_9413);
  not g18672 (n_9414, n9899);
  and g18673 (n9900, n556, n_9414);
  not g18674 (n_9415, n9900);
  and g18675 (n9901, n560, n_9415);
  not g18676 (n_9416, n9901);
  and g18677 (n9902, n564, n_9416);
  not g18678 (n_9417, n9902);
  and g18679 (n9903, n568, n_9417);
  not g18680 (n_9418, n9903);
  and g18681 (n9904, n572, n_9418);
  not g18682 (n_9419, n9904);
  and g18683 (n9905, n576, n_9419);
  not g18684 (n_9420, n9905);
  and g18685 (n9906, n580, n_9420);
  not g18686 (n_9421, n9906);
  and g18687 (n9907, n584, n_9421);
  not g18688 (n_9422, n9907);
  and g18689 (n9908, n588, n_9422);
  not g18690 (n_9423, n9908);
  and g18691 (n9909, n592, n_9423);
  not g18692 (n_9424, n9909);
  and g18693 (n9910, n596, n_9424);
  not g18694 (n_9425, n9910);
  and g18695 (n9911, n600, n_9425);
  not g18696 (n_9426, n9911);
  and g18697 (n9912, n604, n_9426);
  not g18698 (n_9427, n9912);
  and g18699 (n9913, n608, n_9427);
  not g18700 (n_9428, n9913);
  and g18701 (n9914, n612, n_9428);
  not g18702 (n_9429, n9914);
  and g18703 (n9915, n616, n_9429);
  not g18704 (n_9430, n9915);
  and g18705 (n9916, n620, n_9430);
  not g18706 (n_9431, n9916);
  and g18707 (n9917, n624, n_9431);
  not g18708 (n_9432, n9917);
  and g18709 (n9918, n628, n_9432);
  not g18710 (n_9433, n9918);
  and g18711 (n9919, n632, n_9433);
  not g18712 (n_9434, n9919);
  and g18713 (n9920, n636, n_9434);
  not g18714 (n_9435, n9920);
  and g18715 (n9921, n640, n_9435);
  not g18716 (n_9436, n9921);
  and g18717 (n9922, n644, n_9436);
  not g18718 (n_9437, n9922);
  and g18719 (n9923, n648, n_9437);
  and g18720 (n9924, \req[101] , n_472);
  not g18721 (n_9438, n9923);
  and g18722 (\grant[101] , n_9438, n9924);
  not g18723 (n_9439, n994);
  and g18724 (n9926, n659, n_9439);
  not g18725 (n_9440, n9926);
  and g18726 (n9927, n664, n_9440);
  not g18727 (n_9441, n9927);
  and g18728 (n9928, n668, n_9441);
  not g18729 (n_9442, n9928);
  and g18730 (n9929, n672, n_9442);
  not g18731 (n_9443, n9929);
  and g18732 (n9930, n676, n_9443);
  not g18733 (n_9444, n9930);
  and g18734 (n9931, n680, n_9444);
  not g18735 (n_9445, n9931);
  and g18736 (n9932, n684, n_9445);
  not g18737 (n_9446, n9932);
  and g18738 (n9933, n688, n_9446);
  not g18739 (n_9447, n9933);
  and g18740 (n9934, n692, n_9447);
  not g18741 (n_9448, n9934);
  and g18742 (n9935, n696, n_9448);
  not g18743 (n_9449, n9935);
  and g18744 (n9936, n700, n_9449);
  not g18745 (n_9450, n9936);
  and g18746 (n9937, n704, n_9450);
  not g18747 (n_9451, n9937);
  and g18748 (n9938, n708, n_9451);
  not g18749 (n_9452, n9938);
  and g18750 (n9939, n712, n_9452);
  not g18751 (n_9453, n9939);
  and g18752 (n9940, n716, n_9453);
  not g18753 (n_9454, n9940);
  and g18754 (n9941, n720, n_9454);
  not g18755 (n_9455, n9941);
  and g18756 (n9942, n1484, n_9455);
  not g18757 (n_9456, n9942);
  and g18758 (n9943, n1486, n_9456);
  not g18759 (n_9457, n9943);
  and g18760 (n9944, n1750, n_9457);
  not g18761 (n_9458, n9944);
  and g18762 (n9945, n731, n_9458);
  not g18763 (n_9459, n9945);
  and g18764 (n9946, n735, n_9459);
  not g18765 (n_9460, n9946);
  and g18766 (n9947, n739, n_9460);
  not g18767 (n_9461, n9947);
  and g18768 (n9948, n743, n_9461);
  not g18769 (n_9462, n9948);
  and g18770 (n9949, n747, n_9462);
  not g18771 (n_9463, n9949);
  and g18772 (n9950, n751, n_9463);
  not g18773 (n_9464, n9950);
  and g18774 (n9951, n755, n_9464);
  not g18775 (n_9465, n9951);
  and g18776 (n9952, n759, n_9465);
  not g18777 (n_9466, n9952);
  and g18778 (n9953, n763, n_9466);
  not g18779 (n_9467, n9953);
  and g18780 (n9954, n767, n_9467);
  not g18781 (n_9468, n9954);
  and g18782 (n9955, n771, n_9468);
  not g18783 (n_9469, n9955);
  and g18784 (n9956, n775, n_9469);
  not g18785 (n_9470, n9956);
  and g18786 (n9957, n779, n_9470);
  not g18787 (n_9471, n9957);
  and g18788 (n9958, n783, n_9471);
  not g18789 (n_9472, n9958);
  and g18790 (n9959, n787, n_9472);
  not g18791 (n_9473, n9959);
  and g18792 (n9960, n791, n_9473);
  not g18793 (n_9474, n9960);
  and g18794 (n9961, n795, n_9474);
  not g18795 (n_9475, n9961);
  and g18796 (n9962, n799, n_9475);
  not g18797 (n_9476, n9962);
  and g18798 (n9963, n803, n_9476);
  not g18799 (n_9477, n9963);
  and g18800 (n9964, n807, n_9477);
  not g18801 (n_9478, n9964);
  and g18802 (n9965, n811, n_9478);
  not g18803 (n_9479, n9965);
  and g18804 (n9966, n815, n_9479);
  not g18805 (n_9480, n9966);
  and g18806 (n9967, n819, n_9480);
  not g18807 (n_9481, n9967);
  and g18808 (n9968, n823, n_9481);
  not g18809 (n_9482, n9968);
  and g18810 (n9969, n827, n_9482);
  not g18811 (n_9483, n9969);
  and g18812 (n9970, n831, n_9483);
  not g18813 (n_9484, n9970);
  and g18814 (n9971, n835, n_9484);
  not g18815 (n_9485, n9971);
  and g18816 (n9972, n839, n_9485);
  not g18817 (n_9486, n9972);
  and g18818 (n9973, n843, n_9486);
  not g18819 (n_9487, n9973);
  and g18820 (n9974, n847, n_9487);
  not g18821 (n_9488, n9974);
  and g18822 (n9975, n851, n_9488);
  not g18823 (n_9489, n9975);
  and g18824 (n9976, n855, n_9489);
  not g18825 (n_9490, n9976);
  and g18826 (n9977, n859, n_9490);
  not g18827 (n_9491, n9977);
  and g18828 (n9978, n863, n_9491);
  not g18829 (n_9492, n9978);
  and g18830 (n9979, n867, n_9492);
  not g18831 (n_9493, n9979);
  and g18832 (n9980, n871, n_9493);
  not g18833 (n_9494, n9980);
  and g18834 (n9981, n875, n_9494);
  not g18835 (n_9495, n9981);
  and g18836 (n9982, n879, n_9495);
  not g18837 (n_9496, n9982);
  and g18838 (n9983, n883, n_9496);
  not g18839 (n_9497, n9983);
  and g18840 (n9984, n887, n_9497);
  not g18841 (n_9498, n9984);
  and g18842 (n9985, n891, n_9498);
  not g18843 (n_9499, n9985);
  and g18844 (n9986, n895, n_9499);
  not g18845 (n_9500, n9986);
  and g18846 (n9987, n899, n_9500);
  not g18847 (n_9501, n9987);
  and g18848 (n9988, n903, n_9501);
  not g18849 (n_9502, n9988);
  and g18850 (n9989, n907, n_9502);
  not g18851 (n_9503, n9989);
  and g18852 (n9990, n911, n_9503);
  not g18853 (n_9504, n9990);
  and g18854 (n9991, n915, n_9504);
  not g18855 (n_9505, n9991);
  and g18856 (n9992, n919, n_9505);
  not g18857 (n_9506, n9992);
  and g18858 (n9993, n923, n_9506);
  not g18859 (n_9507, n9993);
  and g18860 (n9994, n927, n_9507);
  not g18861 (n_9508, n9994);
  and g18862 (n9995, n931, n_9508);
  not g18863 (n_9509, n9995);
  and g18864 (n9996, n935, n_9509);
  not g18865 (n_9510, n9996);
  and g18866 (n9997, n939, n_9510);
  not g18867 (n_9511, n9997);
  and g18868 (n9998, n943, n_9511);
  not g18869 (n_9512, n9998);
  and g18870 (n9999, n947, n_9512);
  not g18871 (n_9513, n9999);
  and g18872 (n10000, n951, n_9513);
  not g18873 (n_9514, n10000);
  and g18874 (n10001, n955, n_9514);
  not g18875 (n_9515, n10001);
  and g18876 (n10002, n959, n_9515);
  not g18877 (n_9516, n10002);
  and g18878 (n10003, n963, n_9516);
  not g18879 (n_9517, n10003);
  and g18880 (n10004, n967, n_9517);
  not g18881 (n_9518, n10004);
  and g18882 (n10005, n971, n_9518);
  not g18883 (n_9519, n10005);
  and g18884 (n10006, n975, n_9519);
  not g18885 (n_9520, n10006);
  and g18886 (n10007, n979, n_9520);
  not g18887 (n_9521, n10007);
  and g18888 (n10008, n983, n_9521);
  not g18889 (n_9522, n10008);
  and g18890 (n10009, n987, n_9522);
  and g18891 (n10010, \req[102] , n_797);
  not g18892 (n_9523, n10009);
  and g18893 (\grant[102] , n_9523, n10010);
  not g18894 (n_9524, n1331);
  and g18895 (n10012, n998, n_9524);
  not g18896 (n_9525, n10012);
  and g18897 (n10013, n1003, n_9525);
  not g18898 (n_9526, n10013);
  and g18899 (n10014, n1007, n_9526);
  not g18900 (n_9527, n10014);
  and g18901 (n10015, n1011, n_9527);
  not g18902 (n_9528, n10015);
  and g18903 (n10016, n1015, n_9528);
  not g18904 (n_9529, n10016);
  and g18905 (n10017, n1019, n_9529);
  not g18906 (n_9530, n10017);
  and g18907 (n10018, n1023, n_9530);
  not g18908 (n_9531, n10018);
  and g18909 (n10019, n1027, n_9531);
  not g18910 (n_9532, n10019);
  and g18911 (n10020, n1031, n_9532);
  not g18912 (n_9533, n10020);
  and g18913 (n10021, n1035, n_9533);
  not g18914 (n_9534, n10021);
  and g18915 (n10022, n1039, n_9534);
  not g18916 (n_9535, n10022);
  and g18917 (n10023, n1043, n_9535);
  not g18918 (n_9536, n10023);
  and g18919 (n10024, n1047, n_9536);
  not g18920 (n_9537, n10024);
  and g18921 (n10025, n1051, n_9537);
  not g18922 (n_9538, n10025);
  and g18923 (n10026, n1055, n_9538);
  not g18924 (n_9539, n10026);
  and g18925 (n10027, n1059, n_9539);
  not g18926 (n_9540, n10027);
  and g18927 (n10028, n1574, n_9540);
  not g18928 (n_9541, n10028);
  and g18929 (n10029, n1576, n_9541);
  not g18930 (n_9542, n10029);
  and g18931 (n10030, n1837, n_9542);
  not g18932 (n_9543, n10030);
  and g18933 (n10031, n1068, n_9543);
  not g18934 (n_9544, n10031);
  and g18935 (n10032, n1072, n_9544);
  not g18936 (n_9545, n10032);
  and g18937 (n10033, n1076, n_9545);
  not g18938 (n_9546, n10033);
  and g18939 (n10034, n1080, n_9546);
  not g18940 (n_9547, n10034);
  and g18941 (n10035, n1084, n_9547);
  not g18942 (n_9548, n10035);
  and g18943 (n10036, n1088, n_9548);
  not g18944 (n_9549, n10036);
  and g18945 (n10037, n1092, n_9549);
  not g18946 (n_9550, n10037);
  and g18947 (n10038, n1096, n_9550);
  not g18948 (n_9551, n10038);
  and g18949 (n10039, n1100, n_9551);
  not g18950 (n_9552, n10039);
  and g18951 (n10040, n1104, n_9552);
  not g18952 (n_9553, n10040);
  and g18953 (n10041, n1108, n_9553);
  not g18954 (n_9554, n10041);
  and g18955 (n10042, n1112, n_9554);
  not g18956 (n_9555, n10042);
  and g18957 (n10043, n1116, n_9555);
  not g18958 (n_9556, n10043);
  and g18959 (n10044, n1120, n_9556);
  not g18960 (n_9557, n10044);
  and g18961 (n10045, n1124, n_9557);
  not g18962 (n_9558, n10045);
  and g18963 (n10046, n1128, n_9558);
  not g18964 (n_9559, n10046);
  and g18965 (n10047, n1132, n_9559);
  not g18966 (n_9560, n10047);
  and g18967 (n10048, n1136, n_9560);
  not g18968 (n_9561, n10048);
  and g18969 (n10049, n1140, n_9561);
  not g18970 (n_9562, n10049);
  and g18971 (n10050, n1144, n_9562);
  not g18972 (n_9563, n10050);
  and g18973 (n10051, n1148, n_9563);
  not g18974 (n_9564, n10051);
  and g18975 (n10052, n1152, n_9564);
  not g18976 (n_9565, n10052);
  and g18977 (n10053, n1156, n_9565);
  not g18978 (n_9566, n10053);
  and g18979 (n10054, n1160, n_9566);
  not g18980 (n_9567, n10054);
  and g18981 (n10055, n1164, n_9567);
  not g18982 (n_9568, n10055);
  and g18983 (n10056, n1168, n_9568);
  not g18984 (n_9569, n10056);
  and g18985 (n10057, n1172, n_9569);
  not g18986 (n_9570, n10057);
  and g18987 (n10058, n1176, n_9570);
  not g18988 (n_9571, n10058);
  and g18989 (n10059, n1180, n_9571);
  not g18990 (n_9572, n10059);
  and g18991 (n10060, n1184, n_9572);
  not g18992 (n_9573, n10060);
  and g18993 (n10061, n1188, n_9573);
  not g18994 (n_9574, n10061);
  and g18995 (n10062, n1192, n_9574);
  not g18996 (n_9575, n10062);
  and g18997 (n10063, n1196, n_9575);
  not g18998 (n_9576, n10063);
  and g18999 (n10064, n1200, n_9576);
  not g19000 (n_9577, n10064);
  and g19001 (n10065, n1204, n_9577);
  not g19002 (n_9578, n10065);
  and g19003 (n10066, n1208, n_9578);
  not g19004 (n_9579, n10066);
  and g19005 (n10067, n1212, n_9579);
  not g19006 (n_9580, n10067);
  and g19007 (n10068, n1216, n_9580);
  not g19008 (n_9581, n10068);
  and g19009 (n10069, n1220, n_9581);
  not g19010 (n_9582, n10069);
  and g19011 (n10070, n1224, n_9582);
  not g19012 (n_9583, n10070);
  and g19013 (n10071, n1228, n_9583);
  not g19014 (n_9584, n10071);
  and g19015 (n10072, n1232, n_9584);
  not g19016 (n_9585, n10072);
  and g19017 (n10073, n1236, n_9585);
  not g19018 (n_9586, n10073);
  and g19019 (n10074, n1240, n_9586);
  not g19020 (n_9587, n10074);
  and g19021 (n10075, n1244, n_9587);
  not g19022 (n_9588, n10075);
  and g19023 (n10076, n1248, n_9588);
  not g19024 (n_9589, n10076);
  and g19025 (n10077, n1252, n_9589);
  not g19026 (n_9590, n10077);
  and g19027 (n10078, n1256, n_9590);
  not g19028 (n_9591, n10078);
  and g19029 (n10079, n1260, n_9591);
  not g19030 (n_9592, n10079);
  and g19031 (n10080, n1264, n_9592);
  not g19032 (n_9593, n10080);
  and g19033 (n10081, n1268, n_9593);
  not g19034 (n_9594, n10081);
  and g19035 (n10082, n1272, n_9594);
  not g19036 (n_9595, n10082);
  and g19037 (n10083, n1276, n_9595);
  not g19038 (n_9596, n10083);
  and g19039 (n10084, n1280, n_9596);
  not g19040 (n_9597, n10084);
  and g19041 (n10085, n1284, n_9597);
  not g19042 (n_9598, n10085);
  and g19043 (n10086, n1288, n_9598);
  not g19044 (n_9599, n10086);
  and g19045 (n10087, n1292, n_9599);
  not g19046 (n_9600, n10087);
  and g19047 (n10088, n1296, n_9600);
  not g19048 (n_9601, n10088);
  and g19049 (n10089, n1300, n_9601);
  not g19050 (n_9602, n10089);
  and g19051 (n10090, n1304, n_9602);
  not g19052 (n_9603, n10090);
  and g19053 (n10091, n1308, n_9603);
  not g19054 (n_9604, n10091);
  and g19055 (n10092, n1312, n_9604);
  not g19056 (n_9605, n10092);
  and g19057 (n10093, n1316, n_9605);
  not g19058 (n_9606, n10093);
  and g19059 (n10094, n1320, n_9606);
  not g19060 (n_9607, n10094);
  and g19061 (n10095, n1324, n_9607);
  and g19062 (n10096, \req[103] , n_983);
  not g19063 (n_9608, n10095);
  and g19064 (\grant[103] , n_9608, n10096);
  not g19065 (n_9609, n663);
  and g19066 (n10098, n_9609, n1335);
  not g19067 (n_9610, n10098);
  and g19068 (n10099, n1340, n_9610);
  not g19069 (n_9611, n10099);
  and g19070 (n10100, n1344, n_9611);
  not g19071 (n_9612, n10100);
  and g19072 (n10101, n1348, n_9612);
  not g19073 (n_9613, n10101);
  and g19074 (n10102, n1352, n_9613);
  not g19075 (n_9614, n10102);
  and g19076 (n10103, n1356, n_9614);
  not g19077 (n_9615, n10103);
  and g19078 (n10104, n1360, n_9615);
  not g19079 (n_9616, n10104);
  and g19080 (n10105, n1364, n_9616);
  not g19081 (n_9617, n10105);
  and g19082 (n10106, n1368, n_9617);
  not g19083 (n_9618, n10106);
  and g19084 (n10107, n1372, n_9618);
  not g19085 (n_9619, n10107);
  and g19086 (n10108, n1376, n_9619);
  not g19087 (n_9620, n10108);
  and g19088 (n10109, n1380, n_9620);
  not g19089 (n_9621, n10109);
  and g19090 (n10110, n1384, n_9621);
  not g19091 (n_9622, n10110);
  and g19092 (n10111, n1388, n_9622);
  not g19093 (n_9623, n10111);
  and g19094 (n10112, n1392, n_9623);
  not g19095 (n_9624, n10112);
  and g19096 (n10113, n1396, n_9624);
  not g19097 (n_9625, n10113);
  and g19098 (n10114, n1663, n_9625);
  not g19099 (n_9626, n10114);
  and g19100 (n10115, n392, n_9626);
  not g19101 (n_9627, n10115);
  and g19102 (n10116, n396, n_9627);
  not g19103 (n_9628, n10116);
  and g19104 (n10117, n400, n_9628);
  not g19105 (n_9629, n10117);
  and g19106 (n10118, n404, n_9629);
  not g19107 (n_9630, n10118);
  and g19108 (n10119, n408, n_9630);
  not g19109 (n_9631, n10119);
  and g19110 (n10120, n412, n_9631);
  not g19111 (n_9632, n10120);
  and g19112 (n10121, n416, n_9632);
  not g19113 (n_9633, n10121);
  and g19114 (n10122, n420, n_9633);
  not g19115 (n_9634, n10122);
  and g19116 (n10123, n424, n_9634);
  not g19117 (n_9635, n10123);
  and g19118 (n10124, n428, n_9635);
  not g19119 (n_9636, n10124);
  and g19120 (n10125, n432, n_9636);
  not g19121 (n_9637, n10125);
  and g19122 (n10126, n436, n_9637);
  not g19123 (n_9638, n10126);
  and g19124 (n10127, n440, n_9638);
  not g19125 (n_9639, n10127);
  and g19126 (n10128, n444, n_9639);
  not g19127 (n_9640, n10128);
  and g19128 (n10129, n448, n_9640);
  not g19129 (n_9641, n10129);
  and g19130 (n10130, n452, n_9641);
  not g19131 (n_9642, n10130);
  and g19132 (n10131, n456, n_9642);
  not g19133 (n_9643, n10131);
  and g19134 (n10132, n460, n_9643);
  not g19135 (n_9644, n10132);
  and g19136 (n10133, n464, n_9644);
  not g19137 (n_9645, n10133);
  and g19138 (n10134, n468, n_9645);
  not g19139 (n_9646, n10134);
  and g19140 (n10135, n472, n_9646);
  not g19141 (n_9647, n10135);
  and g19142 (n10136, n476, n_9647);
  not g19143 (n_9648, n10136);
  and g19144 (n10137, n480, n_9648);
  not g19145 (n_9649, n10137);
  and g19146 (n10138, n484, n_9649);
  not g19147 (n_9650, n10138);
  and g19148 (n10139, n488, n_9650);
  not g19149 (n_9651, n10139);
  and g19150 (n10140, n492, n_9651);
  not g19151 (n_9652, n10140);
  and g19152 (n10141, n496, n_9652);
  not g19153 (n_9653, n10141);
  and g19154 (n10142, n500, n_9653);
  not g19155 (n_9654, n10142);
  and g19156 (n10143, n504, n_9654);
  not g19157 (n_9655, n10143);
  and g19158 (n10144, n508, n_9655);
  not g19159 (n_9656, n10144);
  and g19160 (n10145, n512, n_9656);
  not g19161 (n_9657, n10145);
  and g19162 (n10146, n516, n_9657);
  not g19163 (n_9658, n10146);
  and g19164 (n10147, n520, n_9658);
  not g19165 (n_9659, n10147);
  and g19166 (n10148, n524, n_9659);
  not g19167 (n_9660, n10148);
  and g19168 (n10149, n528, n_9660);
  not g19169 (n_9661, n10149);
  and g19170 (n10150, n532, n_9661);
  not g19171 (n_9662, n10150);
  and g19172 (n10151, n536, n_9662);
  not g19173 (n_9663, n10151);
  and g19174 (n10152, n540, n_9663);
  not g19175 (n_9664, n10152);
  and g19176 (n10153, n544, n_9664);
  not g19177 (n_9665, n10153);
  and g19178 (n10154, n548, n_9665);
  not g19179 (n_9666, n10154);
  and g19180 (n10155, n552, n_9666);
  not g19181 (n_9667, n10155);
  and g19182 (n10156, n556, n_9667);
  not g19183 (n_9668, n10156);
  and g19184 (n10157, n560, n_9668);
  not g19185 (n_9669, n10157);
  and g19186 (n10158, n564, n_9669);
  not g19187 (n_9670, n10158);
  and g19188 (n10159, n568, n_9670);
  not g19189 (n_9671, n10159);
  and g19190 (n10160, n572, n_9671);
  not g19191 (n_9672, n10160);
  and g19192 (n10161, n576, n_9672);
  not g19193 (n_9673, n10161);
  and g19194 (n10162, n580, n_9673);
  not g19195 (n_9674, n10162);
  and g19196 (n10163, n584, n_9674);
  not g19197 (n_9675, n10163);
  and g19198 (n10164, n588, n_9675);
  not g19199 (n_9676, n10164);
  and g19200 (n10165, n592, n_9676);
  not g19201 (n_9677, n10165);
  and g19202 (n10166, n596, n_9677);
  not g19203 (n_9678, n10166);
  and g19204 (n10167, n600, n_9678);
  not g19205 (n_9679, n10167);
  and g19206 (n10168, n604, n_9679);
  not g19207 (n_9680, n10168);
  and g19208 (n10169, n608, n_9680);
  not g19209 (n_9681, n10169);
  and g19210 (n10170, n612, n_9681);
  not g19211 (n_9682, n10170);
  and g19212 (n10171, n616, n_9682);
  not g19213 (n_9683, n10171);
  and g19214 (n10172, n620, n_9683);
  not g19215 (n_9684, n10172);
  and g19216 (n10173, n624, n_9684);
  not g19217 (n_9685, n10173);
  and g19218 (n10174, n628, n_9685);
  not g19219 (n_9686, n10174);
  and g19220 (n10175, n632, n_9686);
  not g19221 (n_9687, n10175);
  and g19222 (n10176, n636, n_9687);
  not g19223 (n_9688, n10176);
  and g19224 (n10177, n640, n_9688);
  not g19225 (n_9689, n10177);
  and g19226 (n10178, n644, n_9689);
  not g19227 (n_9690, n10178);
  and g19228 (n10179, n648, n_9690);
  not g19229 (n_9691, n10179);
  and g19230 (n10180, n652, n_9691);
  not g19231 (n_9692, n10180);
  and g19232 (n10181, n656, n_9692);
  and g19233 (n10182, \req[104] , n_486);
  not g19234 (n_9693, n10181);
  and g19235 (\grant[104] , n_9693, n10182);
  not g19236 (n_9694, n1002);
  and g19237 (n10184, n667, n_9694);
  not g19238 (n_9695, n10184);
  and g19239 (n10185, n672, n_9695);
  not g19240 (n_9696, n10185);
  and g19241 (n10186, n676, n_9696);
  not g19242 (n_9697, n10186);
  and g19243 (n10187, n680, n_9697);
  not g19244 (n_9698, n10187);
  and g19245 (n10188, n684, n_9698);
  not g19246 (n_9699, n10188);
  and g19247 (n10189, n688, n_9699);
  not g19248 (n_9700, n10189);
  and g19249 (n10190, n692, n_9700);
  not g19250 (n_9701, n10190);
  and g19251 (n10191, n696, n_9701);
  not g19252 (n_9702, n10191);
  and g19253 (n10192, n700, n_9702);
  not g19254 (n_9703, n10192);
  and g19255 (n10193, n704, n_9703);
  not g19256 (n_9704, n10193);
  and g19257 (n10194, n708, n_9704);
  not g19258 (n_9705, n10194);
  and g19259 (n10195, n712, n_9705);
  not g19260 (n_9706, n10195);
  and g19261 (n10196, n716, n_9706);
  not g19262 (n_9707, n10196);
  and g19263 (n10197, n720, n_9707);
  not g19264 (n_9708, n10197);
  and g19265 (n10198, n1484, n_9708);
  not g19266 (n_9709, n10198);
  and g19267 (n10199, n1486, n_9709);
  not g19268 (n_9710, n10199);
  and g19269 (n10200, n1750, n_9710);
  not g19270 (n_9711, n10200);
  and g19271 (n10201, n731, n_9711);
  not g19272 (n_9712, n10201);
  and g19273 (n10202, n735, n_9712);
  not g19274 (n_9713, n10202);
  and g19275 (n10203, n739, n_9713);
  not g19276 (n_9714, n10203);
  and g19277 (n10204, n743, n_9714);
  not g19278 (n_9715, n10204);
  and g19279 (n10205, n747, n_9715);
  not g19280 (n_9716, n10205);
  and g19281 (n10206, n751, n_9716);
  not g19282 (n_9717, n10206);
  and g19283 (n10207, n755, n_9717);
  not g19284 (n_9718, n10207);
  and g19285 (n10208, n759, n_9718);
  not g19286 (n_9719, n10208);
  and g19287 (n10209, n763, n_9719);
  not g19288 (n_9720, n10209);
  and g19289 (n10210, n767, n_9720);
  not g19290 (n_9721, n10210);
  and g19291 (n10211, n771, n_9721);
  not g19292 (n_9722, n10211);
  and g19293 (n10212, n775, n_9722);
  not g19294 (n_9723, n10212);
  and g19295 (n10213, n779, n_9723);
  not g19296 (n_9724, n10213);
  and g19297 (n10214, n783, n_9724);
  not g19298 (n_9725, n10214);
  and g19299 (n10215, n787, n_9725);
  not g19300 (n_9726, n10215);
  and g19301 (n10216, n791, n_9726);
  not g19302 (n_9727, n10216);
  and g19303 (n10217, n795, n_9727);
  not g19304 (n_9728, n10217);
  and g19305 (n10218, n799, n_9728);
  not g19306 (n_9729, n10218);
  and g19307 (n10219, n803, n_9729);
  not g19308 (n_9730, n10219);
  and g19309 (n10220, n807, n_9730);
  not g19310 (n_9731, n10220);
  and g19311 (n10221, n811, n_9731);
  not g19312 (n_9732, n10221);
  and g19313 (n10222, n815, n_9732);
  not g19314 (n_9733, n10222);
  and g19315 (n10223, n819, n_9733);
  not g19316 (n_9734, n10223);
  and g19317 (n10224, n823, n_9734);
  not g19318 (n_9735, n10224);
  and g19319 (n10225, n827, n_9735);
  not g19320 (n_9736, n10225);
  and g19321 (n10226, n831, n_9736);
  not g19322 (n_9737, n10226);
  and g19323 (n10227, n835, n_9737);
  not g19324 (n_9738, n10227);
  and g19325 (n10228, n839, n_9738);
  not g19326 (n_9739, n10228);
  and g19327 (n10229, n843, n_9739);
  not g19328 (n_9740, n10229);
  and g19329 (n10230, n847, n_9740);
  not g19330 (n_9741, n10230);
  and g19331 (n10231, n851, n_9741);
  not g19332 (n_9742, n10231);
  and g19333 (n10232, n855, n_9742);
  not g19334 (n_9743, n10232);
  and g19335 (n10233, n859, n_9743);
  not g19336 (n_9744, n10233);
  and g19337 (n10234, n863, n_9744);
  not g19338 (n_9745, n10234);
  and g19339 (n10235, n867, n_9745);
  not g19340 (n_9746, n10235);
  and g19341 (n10236, n871, n_9746);
  not g19342 (n_9747, n10236);
  and g19343 (n10237, n875, n_9747);
  not g19344 (n_9748, n10237);
  and g19345 (n10238, n879, n_9748);
  not g19346 (n_9749, n10238);
  and g19347 (n10239, n883, n_9749);
  not g19348 (n_9750, n10239);
  and g19349 (n10240, n887, n_9750);
  not g19350 (n_9751, n10240);
  and g19351 (n10241, n891, n_9751);
  not g19352 (n_9752, n10241);
  and g19353 (n10242, n895, n_9752);
  not g19354 (n_9753, n10242);
  and g19355 (n10243, n899, n_9753);
  not g19356 (n_9754, n10243);
  and g19357 (n10244, n903, n_9754);
  not g19358 (n_9755, n10244);
  and g19359 (n10245, n907, n_9755);
  not g19360 (n_9756, n10245);
  and g19361 (n10246, n911, n_9756);
  not g19362 (n_9757, n10246);
  and g19363 (n10247, n915, n_9757);
  not g19364 (n_9758, n10247);
  and g19365 (n10248, n919, n_9758);
  not g19366 (n_9759, n10248);
  and g19367 (n10249, n923, n_9759);
  not g19368 (n_9760, n10249);
  and g19369 (n10250, n927, n_9760);
  not g19370 (n_9761, n10250);
  and g19371 (n10251, n931, n_9761);
  not g19372 (n_9762, n10251);
  and g19373 (n10252, n935, n_9762);
  not g19374 (n_9763, n10252);
  and g19375 (n10253, n939, n_9763);
  not g19376 (n_9764, n10253);
  and g19377 (n10254, n943, n_9764);
  not g19378 (n_9765, n10254);
  and g19379 (n10255, n947, n_9765);
  not g19380 (n_9766, n10255);
  and g19381 (n10256, n951, n_9766);
  not g19382 (n_9767, n10256);
  and g19383 (n10257, n955, n_9767);
  not g19384 (n_9768, n10257);
  and g19385 (n10258, n959, n_9768);
  not g19386 (n_9769, n10258);
  and g19387 (n10259, n963, n_9769);
  not g19388 (n_9770, n10259);
  and g19389 (n10260, n967, n_9770);
  not g19390 (n_9771, n10260);
  and g19391 (n10261, n971, n_9771);
  not g19392 (n_9772, n10261);
  and g19393 (n10262, n975, n_9772);
  not g19394 (n_9773, n10262);
  and g19395 (n10263, n979, n_9773);
  not g19396 (n_9774, n10263);
  and g19397 (n10264, n983, n_9774);
  not g19398 (n_9775, n10264);
  and g19399 (n10265, n987, n_9775);
  not g19400 (n_9776, n10265);
  and g19401 (n10266, n991, n_9776);
  not g19402 (n_9777, n10266);
  and g19403 (n10267, n995, n_9777);
  and g19404 (n10268, \req[105] , n_803);
  not g19405 (n_9778, n10267);
  and g19406 (\grant[105] , n_9778, n10268);
  not g19407 (n_9779, n1339);
  and g19408 (n10270, n1006, n_9779);
  not g19409 (n_9780, n10270);
  and g19410 (n10271, n1011, n_9780);
  not g19411 (n_9781, n10271);
  and g19412 (n10272, n1015, n_9781);
  not g19413 (n_9782, n10272);
  and g19414 (n10273, n1019, n_9782);
  not g19415 (n_9783, n10273);
  and g19416 (n10274, n1023, n_9783);
  not g19417 (n_9784, n10274);
  and g19418 (n10275, n1027, n_9784);
  not g19419 (n_9785, n10275);
  and g19420 (n10276, n1031, n_9785);
  not g19421 (n_9786, n10276);
  and g19422 (n10277, n1035, n_9786);
  not g19423 (n_9787, n10277);
  and g19424 (n10278, n1039, n_9787);
  not g19425 (n_9788, n10278);
  and g19426 (n10279, n1043, n_9788);
  not g19427 (n_9789, n10279);
  and g19428 (n10280, n1047, n_9789);
  not g19429 (n_9790, n10280);
  and g19430 (n10281, n1051, n_9790);
  not g19431 (n_9791, n10281);
  and g19432 (n10282, n1055, n_9791);
  not g19433 (n_9792, n10282);
  and g19434 (n10283, n1059, n_9792);
  not g19435 (n_9793, n10283);
  and g19436 (n10284, n1574, n_9793);
  not g19437 (n_9794, n10284);
  and g19438 (n10285, n1576, n_9794);
  not g19439 (n_9795, n10285);
  and g19440 (n10286, n1837, n_9795);
  not g19441 (n_9796, n10286);
  and g19442 (n10287, n1068, n_9796);
  not g19443 (n_9797, n10287);
  and g19444 (n10288, n1072, n_9797);
  not g19445 (n_9798, n10288);
  and g19446 (n10289, n1076, n_9798);
  not g19447 (n_9799, n10289);
  and g19448 (n10290, n1080, n_9799);
  not g19449 (n_9800, n10290);
  and g19450 (n10291, n1084, n_9800);
  not g19451 (n_9801, n10291);
  and g19452 (n10292, n1088, n_9801);
  not g19453 (n_9802, n10292);
  and g19454 (n10293, n1092, n_9802);
  not g19455 (n_9803, n10293);
  and g19456 (n10294, n1096, n_9803);
  not g19457 (n_9804, n10294);
  and g19458 (n10295, n1100, n_9804);
  not g19459 (n_9805, n10295);
  and g19460 (n10296, n1104, n_9805);
  not g19461 (n_9806, n10296);
  and g19462 (n10297, n1108, n_9806);
  not g19463 (n_9807, n10297);
  and g19464 (n10298, n1112, n_9807);
  not g19465 (n_9808, n10298);
  and g19466 (n10299, n1116, n_9808);
  not g19467 (n_9809, n10299);
  and g19468 (n10300, n1120, n_9809);
  not g19469 (n_9810, n10300);
  and g19470 (n10301, n1124, n_9810);
  not g19471 (n_9811, n10301);
  and g19472 (n10302, n1128, n_9811);
  not g19473 (n_9812, n10302);
  and g19474 (n10303, n1132, n_9812);
  not g19475 (n_9813, n10303);
  and g19476 (n10304, n1136, n_9813);
  not g19477 (n_9814, n10304);
  and g19478 (n10305, n1140, n_9814);
  not g19479 (n_9815, n10305);
  and g19480 (n10306, n1144, n_9815);
  not g19481 (n_9816, n10306);
  and g19482 (n10307, n1148, n_9816);
  not g19483 (n_9817, n10307);
  and g19484 (n10308, n1152, n_9817);
  not g19485 (n_9818, n10308);
  and g19486 (n10309, n1156, n_9818);
  not g19487 (n_9819, n10309);
  and g19488 (n10310, n1160, n_9819);
  not g19489 (n_9820, n10310);
  and g19490 (n10311, n1164, n_9820);
  not g19491 (n_9821, n10311);
  and g19492 (n10312, n1168, n_9821);
  not g19493 (n_9822, n10312);
  and g19494 (n10313, n1172, n_9822);
  not g19495 (n_9823, n10313);
  and g19496 (n10314, n1176, n_9823);
  not g19497 (n_9824, n10314);
  and g19498 (n10315, n1180, n_9824);
  not g19499 (n_9825, n10315);
  and g19500 (n10316, n1184, n_9825);
  not g19501 (n_9826, n10316);
  and g19502 (n10317, n1188, n_9826);
  not g19503 (n_9827, n10317);
  and g19504 (n10318, n1192, n_9827);
  not g19505 (n_9828, n10318);
  and g19506 (n10319, n1196, n_9828);
  not g19507 (n_9829, n10319);
  and g19508 (n10320, n1200, n_9829);
  not g19509 (n_9830, n10320);
  and g19510 (n10321, n1204, n_9830);
  not g19511 (n_9831, n10321);
  and g19512 (n10322, n1208, n_9831);
  not g19513 (n_9832, n10322);
  and g19514 (n10323, n1212, n_9832);
  not g19515 (n_9833, n10323);
  and g19516 (n10324, n1216, n_9833);
  not g19517 (n_9834, n10324);
  and g19518 (n10325, n1220, n_9834);
  not g19519 (n_9835, n10325);
  and g19520 (n10326, n1224, n_9835);
  not g19521 (n_9836, n10326);
  and g19522 (n10327, n1228, n_9836);
  not g19523 (n_9837, n10327);
  and g19524 (n10328, n1232, n_9837);
  not g19525 (n_9838, n10328);
  and g19526 (n10329, n1236, n_9838);
  not g19527 (n_9839, n10329);
  and g19528 (n10330, n1240, n_9839);
  not g19529 (n_9840, n10330);
  and g19530 (n10331, n1244, n_9840);
  not g19531 (n_9841, n10331);
  and g19532 (n10332, n1248, n_9841);
  not g19533 (n_9842, n10332);
  and g19534 (n10333, n1252, n_9842);
  not g19535 (n_9843, n10333);
  and g19536 (n10334, n1256, n_9843);
  not g19537 (n_9844, n10334);
  and g19538 (n10335, n1260, n_9844);
  not g19539 (n_9845, n10335);
  and g19540 (n10336, n1264, n_9845);
  not g19541 (n_9846, n10336);
  and g19542 (n10337, n1268, n_9846);
  not g19543 (n_9847, n10337);
  and g19544 (n10338, n1272, n_9847);
  not g19545 (n_9848, n10338);
  and g19546 (n10339, n1276, n_9848);
  not g19547 (n_9849, n10339);
  and g19548 (n10340, n1280, n_9849);
  not g19549 (n_9850, n10340);
  and g19550 (n10341, n1284, n_9850);
  not g19551 (n_9851, n10341);
  and g19552 (n10342, n1288, n_9851);
  not g19553 (n_9852, n10342);
  and g19554 (n10343, n1292, n_9852);
  not g19555 (n_9853, n10343);
  and g19556 (n10344, n1296, n_9853);
  not g19557 (n_9854, n10344);
  and g19558 (n10345, n1300, n_9854);
  not g19559 (n_9855, n10345);
  and g19560 (n10346, n1304, n_9855);
  not g19561 (n_9856, n10346);
  and g19562 (n10347, n1308, n_9856);
  not g19563 (n_9857, n10347);
  and g19564 (n10348, n1312, n_9857);
  not g19565 (n_9858, n10348);
  and g19566 (n10349, n1316, n_9858);
  not g19567 (n_9859, n10349);
  and g19568 (n10350, n1320, n_9859);
  not g19569 (n_9860, n10350);
  and g19570 (n10351, n1324, n_9860);
  not g19571 (n_9861, n10351);
  and g19572 (n10352, n1328, n_9861);
  not g19573 (n_9862, n10352);
  and g19574 (n10353, n1332, n_9862);
  and g19575 (n10354, \req[106] , n_987);
  not g19576 (n_9863, n10353);
  and g19577 (\grant[106] , n_9863, n10354);
  not g19578 (n_9864, n671);
  and g19579 (n10356, n_9864, n1343);
  not g19580 (n_9865, n10356);
  and g19581 (n10357, n1348, n_9865);
  not g19582 (n_9866, n10357);
  and g19583 (n10358, n1352, n_9866);
  not g19584 (n_9867, n10358);
  and g19585 (n10359, n1356, n_9867);
  not g19586 (n_9868, n10359);
  and g19587 (n10360, n1360, n_9868);
  not g19588 (n_9869, n10360);
  and g19589 (n10361, n1364, n_9869);
  not g19590 (n_9870, n10361);
  and g19591 (n10362, n1368, n_9870);
  not g19592 (n_9871, n10362);
  and g19593 (n10363, n1372, n_9871);
  not g19594 (n_9872, n10363);
  and g19595 (n10364, n1376, n_9872);
  not g19596 (n_9873, n10364);
  and g19597 (n10365, n1380, n_9873);
  not g19598 (n_9874, n10365);
  and g19599 (n10366, n1384, n_9874);
  not g19600 (n_9875, n10366);
  and g19601 (n10367, n1388, n_9875);
  not g19602 (n_9876, n10367);
  and g19603 (n10368, n1392, n_9876);
  not g19604 (n_9877, n10368);
  and g19605 (n10369, n1396, n_9877);
  not g19606 (n_9878, n10369);
  and g19607 (n10370, n1663, n_9878);
  not g19608 (n_9879, n10370);
  and g19609 (n10371, n392, n_9879);
  not g19610 (n_9880, n10371);
  and g19611 (n10372, n396, n_9880);
  not g19612 (n_9881, n10372);
  and g19613 (n10373, n400, n_9881);
  not g19614 (n_9882, n10373);
  and g19615 (n10374, n404, n_9882);
  not g19616 (n_9883, n10374);
  and g19617 (n10375, n408, n_9883);
  not g19618 (n_9884, n10375);
  and g19619 (n10376, n412, n_9884);
  not g19620 (n_9885, n10376);
  and g19621 (n10377, n416, n_9885);
  not g19622 (n_9886, n10377);
  and g19623 (n10378, n420, n_9886);
  not g19624 (n_9887, n10378);
  and g19625 (n10379, n424, n_9887);
  not g19626 (n_9888, n10379);
  and g19627 (n10380, n428, n_9888);
  not g19628 (n_9889, n10380);
  and g19629 (n10381, n432, n_9889);
  not g19630 (n_9890, n10381);
  and g19631 (n10382, n436, n_9890);
  not g19632 (n_9891, n10382);
  and g19633 (n10383, n440, n_9891);
  not g19634 (n_9892, n10383);
  and g19635 (n10384, n444, n_9892);
  not g19636 (n_9893, n10384);
  and g19637 (n10385, n448, n_9893);
  not g19638 (n_9894, n10385);
  and g19639 (n10386, n452, n_9894);
  not g19640 (n_9895, n10386);
  and g19641 (n10387, n456, n_9895);
  not g19642 (n_9896, n10387);
  and g19643 (n10388, n460, n_9896);
  not g19644 (n_9897, n10388);
  and g19645 (n10389, n464, n_9897);
  not g19646 (n_9898, n10389);
  and g19647 (n10390, n468, n_9898);
  not g19648 (n_9899, n10390);
  and g19649 (n10391, n472, n_9899);
  not g19650 (n_9900, n10391);
  and g19651 (n10392, n476, n_9900);
  not g19652 (n_9901, n10392);
  and g19653 (n10393, n480, n_9901);
  not g19654 (n_9902, n10393);
  and g19655 (n10394, n484, n_9902);
  not g19656 (n_9903, n10394);
  and g19657 (n10395, n488, n_9903);
  not g19658 (n_9904, n10395);
  and g19659 (n10396, n492, n_9904);
  not g19660 (n_9905, n10396);
  and g19661 (n10397, n496, n_9905);
  not g19662 (n_9906, n10397);
  and g19663 (n10398, n500, n_9906);
  not g19664 (n_9907, n10398);
  and g19665 (n10399, n504, n_9907);
  not g19666 (n_9908, n10399);
  and g19667 (n10400, n508, n_9908);
  not g19668 (n_9909, n10400);
  and g19669 (n10401, n512, n_9909);
  not g19670 (n_9910, n10401);
  and g19671 (n10402, n516, n_9910);
  not g19672 (n_9911, n10402);
  and g19673 (n10403, n520, n_9911);
  not g19674 (n_9912, n10403);
  and g19675 (n10404, n524, n_9912);
  not g19676 (n_9913, n10404);
  and g19677 (n10405, n528, n_9913);
  not g19678 (n_9914, n10405);
  and g19679 (n10406, n532, n_9914);
  not g19680 (n_9915, n10406);
  and g19681 (n10407, n536, n_9915);
  not g19682 (n_9916, n10407);
  and g19683 (n10408, n540, n_9916);
  not g19684 (n_9917, n10408);
  and g19685 (n10409, n544, n_9917);
  not g19686 (n_9918, n10409);
  and g19687 (n10410, n548, n_9918);
  not g19688 (n_9919, n10410);
  and g19689 (n10411, n552, n_9919);
  not g19690 (n_9920, n10411);
  and g19691 (n10412, n556, n_9920);
  not g19692 (n_9921, n10412);
  and g19693 (n10413, n560, n_9921);
  not g19694 (n_9922, n10413);
  and g19695 (n10414, n564, n_9922);
  not g19696 (n_9923, n10414);
  and g19697 (n10415, n568, n_9923);
  not g19698 (n_9924, n10415);
  and g19699 (n10416, n572, n_9924);
  not g19700 (n_9925, n10416);
  and g19701 (n10417, n576, n_9925);
  not g19702 (n_9926, n10417);
  and g19703 (n10418, n580, n_9926);
  not g19704 (n_9927, n10418);
  and g19705 (n10419, n584, n_9927);
  not g19706 (n_9928, n10419);
  and g19707 (n10420, n588, n_9928);
  not g19708 (n_9929, n10420);
  and g19709 (n10421, n592, n_9929);
  not g19710 (n_9930, n10421);
  and g19711 (n10422, n596, n_9930);
  not g19712 (n_9931, n10422);
  and g19713 (n10423, n600, n_9931);
  not g19714 (n_9932, n10423);
  and g19715 (n10424, n604, n_9932);
  not g19716 (n_9933, n10424);
  and g19717 (n10425, n608, n_9933);
  not g19718 (n_9934, n10425);
  and g19719 (n10426, n612, n_9934);
  not g19720 (n_9935, n10426);
  and g19721 (n10427, n616, n_9935);
  not g19722 (n_9936, n10427);
  and g19723 (n10428, n620, n_9936);
  not g19724 (n_9937, n10428);
  and g19725 (n10429, n624, n_9937);
  not g19726 (n_9938, n10429);
  and g19727 (n10430, n628, n_9938);
  not g19728 (n_9939, n10430);
  and g19729 (n10431, n632, n_9939);
  not g19730 (n_9940, n10431);
  and g19731 (n10432, n636, n_9940);
  not g19732 (n_9941, n10432);
  and g19733 (n10433, n640, n_9941);
  not g19734 (n_9942, n10433);
  and g19735 (n10434, n644, n_9942);
  not g19736 (n_9943, n10434);
  and g19737 (n10435, n648, n_9943);
  not g19738 (n_9944, n10435);
  and g19739 (n10436, n652, n_9944);
  not g19740 (n_9945, n10436);
  and g19741 (n10437, n656, n_9945);
  not g19742 (n_9946, n10437);
  and g19743 (n10438, n660, n_9946);
  not g19744 (n_9947, n10438);
  and g19745 (n10439, n664, n_9947);
  and g19746 (n10440, \req[107] , n_500);
  not g19747 (n_9948, n10439);
  and g19748 (\grant[107] , n_9948, n10440);
  not g19749 (n_9949, n1010);
  and g19750 (n10442, n675, n_9949);
  not g19751 (n_9950, n10442);
  and g19752 (n10443, n680, n_9950);
  not g19753 (n_9951, n10443);
  and g19754 (n10444, n684, n_9951);
  not g19755 (n_9952, n10444);
  and g19756 (n10445, n688, n_9952);
  not g19757 (n_9953, n10445);
  and g19758 (n10446, n692, n_9953);
  not g19759 (n_9954, n10446);
  and g19760 (n10447, n696, n_9954);
  not g19761 (n_9955, n10447);
  and g19762 (n10448, n700, n_9955);
  not g19763 (n_9956, n10448);
  and g19764 (n10449, n704, n_9956);
  not g19765 (n_9957, n10449);
  and g19766 (n10450, n708, n_9957);
  not g19767 (n_9958, n10450);
  and g19768 (n10451, n712, n_9958);
  not g19769 (n_9959, n10451);
  and g19770 (n10452, n716, n_9959);
  not g19771 (n_9960, n10452);
  and g19772 (n10453, n720, n_9960);
  not g19773 (n_9961, n10453);
  and g19774 (n10454, n1484, n_9961);
  not g19775 (n_9962, n10454);
  and g19776 (n10455, n1486, n_9962);
  not g19777 (n_9963, n10455);
  and g19778 (n10456, n1750, n_9963);
  not g19779 (n_9964, n10456);
  and g19780 (n10457, n731, n_9964);
  not g19781 (n_9965, n10457);
  and g19782 (n10458, n735, n_9965);
  not g19783 (n_9966, n10458);
  and g19784 (n10459, n739, n_9966);
  not g19785 (n_9967, n10459);
  and g19786 (n10460, n743, n_9967);
  not g19787 (n_9968, n10460);
  and g19788 (n10461, n747, n_9968);
  not g19789 (n_9969, n10461);
  and g19790 (n10462, n751, n_9969);
  not g19791 (n_9970, n10462);
  and g19792 (n10463, n755, n_9970);
  not g19793 (n_9971, n10463);
  and g19794 (n10464, n759, n_9971);
  not g19795 (n_9972, n10464);
  and g19796 (n10465, n763, n_9972);
  not g19797 (n_9973, n10465);
  and g19798 (n10466, n767, n_9973);
  not g19799 (n_9974, n10466);
  and g19800 (n10467, n771, n_9974);
  not g19801 (n_9975, n10467);
  and g19802 (n10468, n775, n_9975);
  not g19803 (n_9976, n10468);
  and g19804 (n10469, n779, n_9976);
  not g19805 (n_9977, n10469);
  and g19806 (n10470, n783, n_9977);
  not g19807 (n_9978, n10470);
  and g19808 (n10471, n787, n_9978);
  not g19809 (n_9979, n10471);
  and g19810 (n10472, n791, n_9979);
  not g19811 (n_9980, n10472);
  and g19812 (n10473, n795, n_9980);
  not g19813 (n_9981, n10473);
  and g19814 (n10474, n799, n_9981);
  not g19815 (n_9982, n10474);
  and g19816 (n10475, n803, n_9982);
  not g19817 (n_9983, n10475);
  and g19818 (n10476, n807, n_9983);
  not g19819 (n_9984, n10476);
  and g19820 (n10477, n811, n_9984);
  not g19821 (n_9985, n10477);
  and g19822 (n10478, n815, n_9985);
  not g19823 (n_9986, n10478);
  and g19824 (n10479, n819, n_9986);
  not g19825 (n_9987, n10479);
  and g19826 (n10480, n823, n_9987);
  not g19827 (n_9988, n10480);
  and g19828 (n10481, n827, n_9988);
  not g19829 (n_9989, n10481);
  and g19830 (n10482, n831, n_9989);
  not g19831 (n_9990, n10482);
  and g19832 (n10483, n835, n_9990);
  not g19833 (n_9991, n10483);
  and g19834 (n10484, n839, n_9991);
  not g19835 (n_9992, n10484);
  and g19836 (n10485, n843, n_9992);
  not g19837 (n_9993, n10485);
  and g19838 (n10486, n847, n_9993);
  not g19839 (n_9994, n10486);
  and g19840 (n10487, n851, n_9994);
  not g19841 (n_9995, n10487);
  and g19842 (n10488, n855, n_9995);
  not g19843 (n_9996, n10488);
  and g19844 (n10489, n859, n_9996);
  not g19845 (n_9997, n10489);
  and g19846 (n10490, n863, n_9997);
  not g19847 (n_9998, n10490);
  and g19848 (n10491, n867, n_9998);
  not g19849 (n_9999, n10491);
  and g19850 (n10492, n871, n_9999);
  not g19851 (n_10000, n10492);
  and g19852 (n10493, n875, n_10000);
  not g19853 (n_10001, n10493);
  and g19854 (n10494, n879, n_10001);
  not g19855 (n_10002, n10494);
  and g19856 (n10495, n883, n_10002);
  not g19857 (n_10003, n10495);
  and g19858 (n10496, n887, n_10003);
  not g19859 (n_10004, n10496);
  and g19860 (n10497, n891, n_10004);
  not g19861 (n_10005, n10497);
  and g19862 (n10498, n895, n_10005);
  not g19863 (n_10006, n10498);
  and g19864 (n10499, n899, n_10006);
  not g19865 (n_10007, n10499);
  and g19866 (n10500, n903, n_10007);
  not g19867 (n_10008, n10500);
  and g19868 (n10501, n907, n_10008);
  not g19869 (n_10009, n10501);
  and g19870 (n10502, n911, n_10009);
  not g19871 (n_10010, n10502);
  and g19872 (n10503, n915, n_10010);
  not g19873 (n_10011, n10503);
  and g19874 (n10504, n919, n_10011);
  not g19875 (n_10012, n10504);
  and g19876 (n10505, n923, n_10012);
  not g19877 (n_10013, n10505);
  and g19878 (n10506, n927, n_10013);
  not g19879 (n_10014, n10506);
  and g19880 (n10507, n931, n_10014);
  not g19881 (n_10015, n10507);
  and g19882 (n10508, n935, n_10015);
  not g19883 (n_10016, n10508);
  and g19884 (n10509, n939, n_10016);
  not g19885 (n_10017, n10509);
  and g19886 (n10510, n943, n_10017);
  not g19887 (n_10018, n10510);
  and g19888 (n10511, n947, n_10018);
  not g19889 (n_10019, n10511);
  and g19890 (n10512, n951, n_10019);
  not g19891 (n_10020, n10512);
  and g19892 (n10513, n955, n_10020);
  not g19893 (n_10021, n10513);
  and g19894 (n10514, n959, n_10021);
  not g19895 (n_10022, n10514);
  and g19896 (n10515, n963, n_10022);
  not g19897 (n_10023, n10515);
  and g19898 (n10516, n967, n_10023);
  not g19899 (n_10024, n10516);
  and g19900 (n10517, n971, n_10024);
  not g19901 (n_10025, n10517);
  and g19902 (n10518, n975, n_10025);
  not g19903 (n_10026, n10518);
  and g19904 (n10519, n979, n_10026);
  not g19905 (n_10027, n10519);
  and g19906 (n10520, n983, n_10027);
  not g19907 (n_10028, n10520);
  and g19908 (n10521, n987, n_10028);
  not g19909 (n_10029, n10521);
  and g19910 (n10522, n991, n_10029);
  not g19911 (n_10030, n10522);
  and g19912 (n10523, n995, n_10030);
  not g19913 (n_10031, n10523);
  and g19914 (n10524, n999, n_10031);
  not g19915 (n_10032, n10524);
  and g19916 (n10525, n1003, n_10032);
  and g19917 (n10526, \req[108] , n_809);
  not g19918 (n_10033, n10525);
  and g19919 (\grant[108] , n_10033, n10526);
  not g19920 (n_10034, n1347);
  and g19921 (n10528, n1014, n_10034);
  not g19922 (n_10035, n10528);
  and g19923 (n10529, n1019, n_10035);
  not g19924 (n_10036, n10529);
  and g19925 (n10530, n1023, n_10036);
  not g19926 (n_10037, n10530);
  and g19927 (n10531, n1027, n_10037);
  not g19928 (n_10038, n10531);
  and g19929 (n10532, n1031, n_10038);
  not g19930 (n_10039, n10532);
  and g19931 (n10533, n1035, n_10039);
  not g19932 (n_10040, n10533);
  and g19933 (n10534, n1039, n_10040);
  not g19934 (n_10041, n10534);
  and g19935 (n10535, n1043, n_10041);
  not g19936 (n_10042, n10535);
  and g19937 (n10536, n1047, n_10042);
  not g19938 (n_10043, n10536);
  and g19939 (n10537, n1051, n_10043);
  not g19940 (n_10044, n10537);
  and g19941 (n10538, n1055, n_10044);
  not g19942 (n_10045, n10538);
  and g19943 (n10539, n1059, n_10045);
  not g19944 (n_10046, n10539);
  and g19945 (n10540, n1574, n_10046);
  not g19946 (n_10047, n10540);
  and g19947 (n10541, n1576, n_10047);
  not g19948 (n_10048, n10541);
  and g19949 (n10542, n1837, n_10048);
  not g19950 (n_10049, n10542);
  and g19951 (n10543, n1068, n_10049);
  not g19952 (n_10050, n10543);
  and g19953 (n10544, n1072, n_10050);
  not g19954 (n_10051, n10544);
  and g19955 (n10545, n1076, n_10051);
  not g19956 (n_10052, n10545);
  and g19957 (n10546, n1080, n_10052);
  not g19958 (n_10053, n10546);
  and g19959 (n10547, n1084, n_10053);
  not g19960 (n_10054, n10547);
  and g19961 (n10548, n1088, n_10054);
  not g19962 (n_10055, n10548);
  and g19963 (n10549, n1092, n_10055);
  not g19964 (n_10056, n10549);
  and g19965 (n10550, n1096, n_10056);
  not g19966 (n_10057, n10550);
  and g19967 (n10551, n1100, n_10057);
  not g19968 (n_10058, n10551);
  and g19969 (n10552, n1104, n_10058);
  not g19970 (n_10059, n10552);
  and g19971 (n10553, n1108, n_10059);
  not g19972 (n_10060, n10553);
  and g19973 (n10554, n1112, n_10060);
  not g19974 (n_10061, n10554);
  and g19975 (n10555, n1116, n_10061);
  not g19976 (n_10062, n10555);
  and g19977 (n10556, n1120, n_10062);
  not g19978 (n_10063, n10556);
  and g19979 (n10557, n1124, n_10063);
  not g19980 (n_10064, n10557);
  and g19981 (n10558, n1128, n_10064);
  not g19982 (n_10065, n10558);
  and g19983 (n10559, n1132, n_10065);
  not g19984 (n_10066, n10559);
  and g19985 (n10560, n1136, n_10066);
  not g19986 (n_10067, n10560);
  and g19987 (n10561, n1140, n_10067);
  not g19988 (n_10068, n10561);
  and g19989 (n10562, n1144, n_10068);
  not g19990 (n_10069, n10562);
  and g19991 (n10563, n1148, n_10069);
  not g19992 (n_10070, n10563);
  and g19993 (n10564, n1152, n_10070);
  not g19994 (n_10071, n10564);
  and g19995 (n10565, n1156, n_10071);
  not g19996 (n_10072, n10565);
  and g19997 (n10566, n1160, n_10072);
  not g19998 (n_10073, n10566);
  and g19999 (n10567, n1164, n_10073);
  not g20000 (n_10074, n10567);
  and g20001 (n10568, n1168, n_10074);
  not g20002 (n_10075, n10568);
  and g20003 (n10569, n1172, n_10075);
  not g20004 (n_10076, n10569);
  and g20005 (n10570, n1176, n_10076);
  not g20006 (n_10077, n10570);
  and g20007 (n10571, n1180, n_10077);
  not g20008 (n_10078, n10571);
  and g20009 (n10572, n1184, n_10078);
  not g20010 (n_10079, n10572);
  and g20011 (n10573, n1188, n_10079);
  not g20012 (n_10080, n10573);
  and g20013 (n10574, n1192, n_10080);
  not g20014 (n_10081, n10574);
  and g20015 (n10575, n1196, n_10081);
  not g20016 (n_10082, n10575);
  and g20017 (n10576, n1200, n_10082);
  not g20018 (n_10083, n10576);
  and g20019 (n10577, n1204, n_10083);
  not g20020 (n_10084, n10577);
  and g20021 (n10578, n1208, n_10084);
  not g20022 (n_10085, n10578);
  and g20023 (n10579, n1212, n_10085);
  not g20024 (n_10086, n10579);
  and g20025 (n10580, n1216, n_10086);
  not g20026 (n_10087, n10580);
  and g20027 (n10581, n1220, n_10087);
  not g20028 (n_10088, n10581);
  and g20029 (n10582, n1224, n_10088);
  not g20030 (n_10089, n10582);
  and g20031 (n10583, n1228, n_10089);
  not g20032 (n_10090, n10583);
  and g20033 (n10584, n1232, n_10090);
  not g20034 (n_10091, n10584);
  and g20035 (n10585, n1236, n_10091);
  not g20036 (n_10092, n10585);
  and g20037 (n10586, n1240, n_10092);
  not g20038 (n_10093, n10586);
  and g20039 (n10587, n1244, n_10093);
  not g20040 (n_10094, n10587);
  and g20041 (n10588, n1248, n_10094);
  not g20042 (n_10095, n10588);
  and g20043 (n10589, n1252, n_10095);
  not g20044 (n_10096, n10589);
  and g20045 (n10590, n1256, n_10096);
  not g20046 (n_10097, n10590);
  and g20047 (n10591, n1260, n_10097);
  not g20048 (n_10098, n10591);
  and g20049 (n10592, n1264, n_10098);
  not g20050 (n_10099, n10592);
  and g20051 (n10593, n1268, n_10099);
  not g20052 (n_10100, n10593);
  and g20053 (n10594, n1272, n_10100);
  not g20054 (n_10101, n10594);
  and g20055 (n10595, n1276, n_10101);
  not g20056 (n_10102, n10595);
  and g20057 (n10596, n1280, n_10102);
  not g20058 (n_10103, n10596);
  and g20059 (n10597, n1284, n_10103);
  not g20060 (n_10104, n10597);
  and g20061 (n10598, n1288, n_10104);
  not g20062 (n_10105, n10598);
  and g20063 (n10599, n1292, n_10105);
  not g20064 (n_10106, n10599);
  and g20065 (n10600, n1296, n_10106);
  not g20066 (n_10107, n10600);
  and g20067 (n10601, n1300, n_10107);
  not g20068 (n_10108, n10601);
  and g20069 (n10602, n1304, n_10108);
  not g20070 (n_10109, n10602);
  and g20071 (n10603, n1308, n_10109);
  not g20072 (n_10110, n10603);
  and g20073 (n10604, n1312, n_10110);
  not g20074 (n_10111, n10604);
  and g20075 (n10605, n1316, n_10111);
  not g20076 (n_10112, n10605);
  and g20077 (n10606, n1320, n_10112);
  not g20078 (n_10113, n10606);
  and g20079 (n10607, n1324, n_10113);
  not g20080 (n_10114, n10607);
  and g20081 (n10608, n1328, n_10114);
  not g20082 (n_10115, n10608);
  and g20083 (n10609, n1332, n_10115);
  not g20084 (n_10116, n10609);
  and g20085 (n10610, n1336, n_10116);
  not g20086 (n_10117, n10610);
  and g20087 (n10611, n1340, n_10117);
  and g20088 (n10612, \req[109] , n_991);
  not g20089 (n_10118, n10611);
  and g20090 (\grant[109] , n_10118, n10612);
  not g20091 (n_10119, n679);
  and g20092 (n10614, n_10119, n1351);
  not g20093 (n_10120, n10614);
  and g20094 (n10615, n1356, n_10120);
  not g20095 (n_10121, n10615);
  and g20096 (n10616, n1360, n_10121);
  not g20097 (n_10122, n10616);
  and g20098 (n10617, n1364, n_10122);
  not g20099 (n_10123, n10617);
  and g20100 (n10618, n1368, n_10123);
  not g20101 (n_10124, n10618);
  and g20102 (n10619, n1372, n_10124);
  not g20103 (n_10125, n10619);
  and g20104 (n10620, n1376, n_10125);
  not g20105 (n_10126, n10620);
  and g20106 (n10621, n1380, n_10126);
  not g20107 (n_10127, n10621);
  and g20108 (n10622, n1384, n_10127);
  not g20109 (n_10128, n10622);
  and g20110 (n10623, n1388, n_10128);
  not g20111 (n_10129, n10623);
  and g20112 (n10624, n1392, n_10129);
  not g20113 (n_10130, n10624);
  and g20114 (n10625, n1396, n_10130);
  not g20115 (n_10131, n10625);
  and g20116 (n10626, n1663, n_10131);
  not g20117 (n_10132, n10626);
  and g20118 (n10627, n392, n_10132);
  not g20119 (n_10133, n10627);
  and g20120 (n10628, n396, n_10133);
  not g20121 (n_10134, n10628);
  and g20122 (n10629, n400, n_10134);
  not g20123 (n_10135, n10629);
  and g20124 (n10630, n404, n_10135);
  not g20125 (n_10136, n10630);
  and g20126 (n10631, n408, n_10136);
  not g20127 (n_10137, n10631);
  and g20128 (n10632, n412, n_10137);
  not g20129 (n_10138, n10632);
  and g20130 (n10633, n416, n_10138);
  not g20131 (n_10139, n10633);
  and g20132 (n10634, n420, n_10139);
  not g20133 (n_10140, n10634);
  and g20134 (n10635, n424, n_10140);
  not g20135 (n_10141, n10635);
  and g20136 (n10636, n428, n_10141);
  not g20137 (n_10142, n10636);
  and g20138 (n10637, n432, n_10142);
  not g20139 (n_10143, n10637);
  and g20140 (n10638, n436, n_10143);
  not g20141 (n_10144, n10638);
  and g20142 (n10639, n440, n_10144);
  not g20143 (n_10145, n10639);
  and g20144 (n10640, n444, n_10145);
  not g20145 (n_10146, n10640);
  and g20146 (n10641, n448, n_10146);
  not g20147 (n_10147, n10641);
  and g20148 (n10642, n452, n_10147);
  not g20149 (n_10148, n10642);
  and g20150 (n10643, n456, n_10148);
  not g20151 (n_10149, n10643);
  and g20152 (n10644, n460, n_10149);
  not g20153 (n_10150, n10644);
  and g20154 (n10645, n464, n_10150);
  not g20155 (n_10151, n10645);
  and g20156 (n10646, n468, n_10151);
  not g20157 (n_10152, n10646);
  and g20158 (n10647, n472, n_10152);
  not g20159 (n_10153, n10647);
  and g20160 (n10648, n476, n_10153);
  not g20161 (n_10154, n10648);
  and g20162 (n10649, n480, n_10154);
  not g20163 (n_10155, n10649);
  and g20164 (n10650, n484, n_10155);
  not g20165 (n_10156, n10650);
  and g20166 (n10651, n488, n_10156);
  not g20167 (n_10157, n10651);
  and g20168 (n10652, n492, n_10157);
  not g20169 (n_10158, n10652);
  and g20170 (n10653, n496, n_10158);
  not g20171 (n_10159, n10653);
  and g20172 (n10654, n500, n_10159);
  not g20173 (n_10160, n10654);
  and g20174 (n10655, n504, n_10160);
  not g20175 (n_10161, n10655);
  and g20176 (n10656, n508, n_10161);
  not g20177 (n_10162, n10656);
  and g20178 (n10657, n512, n_10162);
  not g20179 (n_10163, n10657);
  and g20180 (n10658, n516, n_10163);
  not g20181 (n_10164, n10658);
  and g20182 (n10659, n520, n_10164);
  not g20183 (n_10165, n10659);
  and g20184 (n10660, n524, n_10165);
  not g20185 (n_10166, n10660);
  and g20186 (n10661, n528, n_10166);
  not g20187 (n_10167, n10661);
  and g20188 (n10662, n532, n_10167);
  not g20189 (n_10168, n10662);
  and g20190 (n10663, n536, n_10168);
  not g20191 (n_10169, n10663);
  and g20192 (n10664, n540, n_10169);
  not g20193 (n_10170, n10664);
  and g20194 (n10665, n544, n_10170);
  not g20195 (n_10171, n10665);
  and g20196 (n10666, n548, n_10171);
  not g20197 (n_10172, n10666);
  and g20198 (n10667, n552, n_10172);
  not g20199 (n_10173, n10667);
  and g20200 (n10668, n556, n_10173);
  not g20201 (n_10174, n10668);
  and g20202 (n10669, n560, n_10174);
  not g20203 (n_10175, n10669);
  and g20204 (n10670, n564, n_10175);
  not g20205 (n_10176, n10670);
  and g20206 (n10671, n568, n_10176);
  not g20207 (n_10177, n10671);
  and g20208 (n10672, n572, n_10177);
  not g20209 (n_10178, n10672);
  and g20210 (n10673, n576, n_10178);
  not g20211 (n_10179, n10673);
  and g20212 (n10674, n580, n_10179);
  not g20213 (n_10180, n10674);
  and g20214 (n10675, n584, n_10180);
  not g20215 (n_10181, n10675);
  and g20216 (n10676, n588, n_10181);
  not g20217 (n_10182, n10676);
  and g20218 (n10677, n592, n_10182);
  not g20219 (n_10183, n10677);
  and g20220 (n10678, n596, n_10183);
  not g20221 (n_10184, n10678);
  and g20222 (n10679, n600, n_10184);
  not g20223 (n_10185, n10679);
  and g20224 (n10680, n604, n_10185);
  not g20225 (n_10186, n10680);
  and g20226 (n10681, n608, n_10186);
  not g20227 (n_10187, n10681);
  and g20228 (n10682, n612, n_10187);
  not g20229 (n_10188, n10682);
  and g20230 (n10683, n616, n_10188);
  not g20231 (n_10189, n10683);
  and g20232 (n10684, n620, n_10189);
  not g20233 (n_10190, n10684);
  and g20234 (n10685, n624, n_10190);
  not g20235 (n_10191, n10685);
  and g20236 (n10686, n628, n_10191);
  not g20237 (n_10192, n10686);
  and g20238 (n10687, n632, n_10192);
  not g20239 (n_10193, n10687);
  and g20240 (n10688, n636, n_10193);
  not g20241 (n_10194, n10688);
  and g20242 (n10689, n640, n_10194);
  not g20243 (n_10195, n10689);
  and g20244 (n10690, n644, n_10195);
  not g20245 (n_10196, n10690);
  and g20246 (n10691, n648, n_10196);
  not g20247 (n_10197, n10691);
  and g20248 (n10692, n652, n_10197);
  not g20249 (n_10198, n10692);
  and g20250 (n10693, n656, n_10198);
  not g20251 (n_10199, n10693);
  and g20252 (n10694, n660, n_10199);
  not g20253 (n_10200, n10694);
  and g20254 (n10695, n664, n_10200);
  not g20255 (n_10201, n10695);
  and g20256 (n10696, n668, n_10201);
  not g20257 (n_10202, n10696);
  and g20258 (n10697, n672, n_10202);
  and g20259 (n10698, \req[110] , n_514);
  not g20260 (n_10203, n10697);
  and g20261 (\grant[110] , n_10203, n10698);
  not g20262 (n_10204, n1018);
  and g20263 (n10700, n683, n_10204);
  not g20264 (n_10205, n10700);
  and g20265 (n10701, n688, n_10205);
  not g20266 (n_10206, n10701);
  and g20267 (n10702, n692, n_10206);
  not g20268 (n_10207, n10702);
  and g20269 (n10703, n696, n_10207);
  not g20270 (n_10208, n10703);
  and g20271 (n10704, n700, n_10208);
  not g20272 (n_10209, n10704);
  and g20273 (n10705, n704, n_10209);
  not g20274 (n_10210, n10705);
  and g20275 (n10706, n708, n_10210);
  not g20276 (n_10211, n10706);
  and g20277 (n10707, n712, n_10211);
  not g20278 (n_10212, n10707);
  and g20279 (n10708, n716, n_10212);
  not g20280 (n_10213, n10708);
  and g20281 (n10709, n720, n_10213);
  not g20282 (n_10214, n10709);
  and g20283 (n10710, n1484, n_10214);
  not g20284 (n_10215, n10710);
  and g20285 (n10711, n1486, n_10215);
  not g20286 (n_10216, n10711);
  and g20287 (n10712, n1750, n_10216);
  not g20288 (n_10217, n10712);
  and g20289 (n10713, n731, n_10217);
  not g20290 (n_10218, n10713);
  and g20291 (n10714, n735, n_10218);
  not g20292 (n_10219, n10714);
  and g20293 (n10715, n739, n_10219);
  not g20294 (n_10220, n10715);
  and g20295 (n10716, n743, n_10220);
  not g20296 (n_10221, n10716);
  and g20297 (n10717, n747, n_10221);
  not g20298 (n_10222, n10717);
  and g20299 (n10718, n751, n_10222);
  not g20300 (n_10223, n10718);
  and g20301 (n10719, n755, n_10223);
  not g20302 (n_10224, n10719);
  and g20303 (n10720, n759, n_10224);
  not g20304 (n_10225, n10720);
  and g20305 (n10721, n763, n_10225);
  not g20306 (n_10226, n10721);
  and g20307 (n10722, n767, n_10226);
  not g20308 (n_10227, n10722);
  and g20309 (n10723, n771, n_10227);
  not g20310 (n_10228, n10723);
  and g20311 (n10724, n775, n_10228);
  not g20312 (n_10229, n10724);
  and g20313 (n10725, n779, n_10229);
  not g20314 (n_10230, n10725);
  and g20315 (n10726, n783, n_10230);
  not g20316 (n_10231, n10726);
  and g20317 (n10727, n787, n_10231);
  not g20318 (n_10232, n10727);
  and g20319 (n10728, n791, n_10232);
  not g20320 (n_10233, n10728);
  and g20321 (n10729, n795, n_10233);
  not g20322 (n_10234, n10729);
  and g20323 (n10730, n799, n_10234);
  not g20324 (n_10235, n10730);
  and g20325 (n10731, n803, n_10235);
  not g20326 (n_10236, n10731);
  and g20327 (n10732, n807, n_10236);
  not g20328 (n_10237, n10732);
  and g20329 (n10733, n811, n_10237);
  not g20330 (n_10238, n10733);
  and g20331 (n10734, n815, n_10238);
  not g20332 (n_10239, n10734);
  and g20333 (n10735, n819, n_10239);
  not g20334 (n_10240, n10735);
  and g20335 (n10736, n823, n_10240);
  not g20336 (n_10241, n10736);
  and g20337 (n10737, n827, n_10241);
  not g20338 (n_10242, n10737);
  and g20339 (n10738, n831, n_10242);
  not g20340 (n_10243, n10738);
  and g20341 (n10739, n835, n_10243);
  not g20342 (n_10244, n10739);
  and g20343 (n10740, n839, n_10244);
  not g20344 (n_10245, n10740);
  and g20345 (n10741, n843, n_10245);
  not g20346 (n_10246, n10741);
  and g20347 (n10742, n847, n_10246);
  not g20348 (n_10247, n10742);
  and g20349 (n10743, n851, n_10247);
  not g20350 (n_10248, n10743);
  and g20351 (n10744, n855, n_10248);
  not g20352 (n_10249, n10744);
  and g20353 (n10745, n859, n_10249);
  not g20354 (n_10250, n10745);
  and g20355 (n10746, n863, n_10250);
  not g20356 (n_10251, n10746);
  and g20357 (n10747, n867, n_10251);
  not g20358 (n_10252, n10747);
  and g20359 (n10748, n871, n_10252);
  not g20360 (n_10253, n10748);
  and g20361 (n10749, n875, n_10253);
  not g20362 (n_10254, n10749);
  and g20363 (n10750, n879, n_10254);
  not g20364 (n_10255, n10750);
  and g20365 (n10751, n883, n_10255);
  not g20366 (n_10256, n10751);
  and g20367 (n10752, n887, n_10256);
  not g20368 (n_10257, n10752);
  and g20369 (n10753, n891, n_10257);
  not g20370 (n_10258, n10753);
  and g20371 (n10754, n895, n_10258);
  not g20372 (n_10259, n10754);
  and g20373 (n10755, n899, n_10259);
  not g20374 (n_10260, n10755);
  and g20375 (n10756, n903, n_10260);
  not g20376 (n_10261, n10756);
  and g20377 (n10757, n907, n_10261);
  not g20378 (n_10262, n10757);
  and g20379 (n10758, n911, n_10262);
  not g20380 (n_10263, n10758);
  and g20381 (n10759, n915, n_10263);
  not g20382 (n_10264, n10759);
  and g20383 (n10760, n919, n_10264);
  not g20384 (n_10265, n10760);
  and g20385 (n10761, n923, n_10265);
  not g20386 (n_10266, n10761);
  and g20387 (n10762, n927, n_10266);
  not g20388 (n_10267, n10762);
  and g20389 (n10763, n931, n_10267);
  not g20390 (n_10268, n10763);
  and g20391 (n10764, n935, n_10268);
  not g20392 (n_10269, n10764);
  and g20393 (n10765, n939, n_10269);
  not g20394 (n_10270, n10765);
  and g20395 (n10766, n943, n_10270);
  not g20396 (n_10271, n10766);
  and g20397 (n10767, n947, n_10271);
  not g20398 (n_10272, n10767);
  and g20399 (n10768, n951, n_10272);
  not g20400 (n_10273, n10768);
  and g20401 (n10769, n955, n_10273);
  not g20402 (n_10274, n10769);
  and g20403 (n10770, n959, n_10274);
  not g20404 (n_10275, n10770);
  and g20405 (n10771, n963, n_10275);
  not g20406 (n_10276, n10771);
  and g20407 (n10772, n967, n_10276);
  not g20408 (n_10277, n10772);
  and g20409 (n10773, n971, n_10277);
  not g20410 (n_10278, n10773);
  and g20411 (n10774, n975, n_10278);
  not g20412 (n_10279, n10774);
  and g20413 (n10775, n979, n_10279);
  not g20414 (n_10280, n10775);
  and g20415 (n10776, n983, n_10280);
  not g20416 (n_10281, n10776);
  and g20417 (n10777, n987, n_10281);
  not g20418 (n_10282, n10777);
  and g20419 (n10778, n991, n_10282);
  not g20420 (n_10283, n10778);
  and g20421 (n10779, n995, n_10283);
  not g20422 (n_10284, n10779);
  and g20423 (n10780, n999, n_10284);
  not g20424 (n_10285, n10780);
  and g20425 (n10781, n1003, n_10285);
  not g20426 (n_10286, n10781);
  and g20427 (n10782, n1007, n_10286);
  not g20428 (n_10287, n10782);
  and g20429 (n10783, n1011, n_10287);
  and g20430 (n10784, \req[111] , n_815);
  not g20431 (n_10288, n10783);
  and g20432 (\grant[111] , n_10288, n10784);
  not g20433 (n_10289, n1355);
  and g20434 (n10786, n1022, n_10289);
  not g20435 (n_10290, n10786);
  and g20436 (n10787, n1027, n_10290);
  not g20437 (n_10291, n10787);
  and g20438 (n10788, n1031, n_10291);
  not g20439 (n_10292, n10788);
  and g20440 (n10789, n1035, n_10292);
  not g20441 (n_10293, n10789);
  and g20442 (n10790, n1039, n_10293);
  not g20443 (n_10294, n10790);
  and g20444 (n10791, n1043, n_10294);
  not g20445 (n_10295, n10791);
  and g20446 (n10792, n1047, n_10295);
  not g20447 (n_10296, n10792);
  and g20448 (n10793, n1051, n_10296);
  not g20449 (n_10297, n10793);
  and g20450 (n10794, n1055, n_10297);
  not g20451 (n_10298, n10794);
  and g20452 (n10795, n1059, n_10298);
  not g20453 (n_10299, n10795);
  and g20454 (n10796, n1574, n_10299);
  not g20455 (n_10300, n10796);
  and g20456 (n10797, n1576, n_10300);
  not g20457 (n_10301, n10797);
  and g20458 (n10798, n1837, n_10301);
  not g20459 (n_10302, n10798);
  and g20460 (n10799, n1068, n_10302);
  not g20461 (n_10303, n10799);
  and g20462 (n10800, n1072, n_10303);
  not g20463 (n_10304, n10800);
  and g20464 (n10801, n1076, n_10304);
  not g20465 (n_10305, n10801);
  and g20466 (n10802, n1080, n_10305);
  not g20467 (n_10306, n10802);
  and g20468 (n10803, n1084, n_10306);
  not g20469 (n_10307, n10803);
  and g20470 (n10804, n1088, n_10307);
  not g20471 (n_10308, n10804);
  and g20472 (n10805, n1092, n_10308);
  not g20473 (n_10309, n10805);
  and g20474 (n10806, n1096, n_10309);
  not g20475 (n_10310, n10806);
  and g20476 (n10807, n1100, n_10310);
  not g20477 (n_10311, n10807);
  and g20478 (n10808, n1104, n_10311);
  not g20479 (n_10312, n10808);
  and g20480 (n10809, n1108, n_10312);
  not g20481 (n_10313, n10809);
  and g20482 (n10810, n1112, n_10313);
  not g20483 (n_10314, n10810);
  and g20484 (n10811, n1116, n_10314);
  not g20485 (n_10315, n10811);
  and g20486 (n10812, n1120, n_10315);
  not g20487 (n_10316, n10812);
  and g20488 (n10813, n1124, n_10316);
  not g20489 (n_10317, n10813);
  and g20490 (n10814, n1128, n_10317);
  not g20491 (n_10318, n10814);
  and g20492 (n10815, n1132, n_10318);
  not g20493 (n_10319, n10815);
  and g20494 (n10816, n1136, n_10319);
  not g20495 (n_10320, n10816);
  and g20496 (n10817, n1140, n_10320);
  not g20497 (n_10321, n10817);
  and g20498 (n10818, n1144, n_10321);
  not g20499 (n_10322, n10818);
  and g20500 (n10819, n1148, n_10322);
  not g20501 (n_10323, n10819);
  and g20502 (n10820, n1152, n_10323);
  not g20503 (n_10324, n10820);
  and g20504 (n10821, n1156, n_10324);
  not g20505 (n_10325, n10821);
  and g20506 (n10822, n1160, n_10325);
  not g20507 (n_10326, n10822);
  and g20508 (n10823, n1164, n_10326);
  not g20509 (n_10327, n10823);
  and g20510 (n10824, n1168, n_10327);
  not g20511 (n_10328, n10824);
  and g20512 (n10825, n1172, n_10328);
  not g20513 (n_10329, n10825);
  and g20514 (n10826, n1176, n_10329);
  not g20515 (n_10330, n10826);
  and g20516 (n10827, n1180, n_10330);
  not g20517 (n_10331, n10827);
  and g20518 (n10828, n1184, n_10331);
  not g20519 (n_10332, n10828);
  and g20520 (n10829, n1188, n_10332);
  not g20521 (n_10333, n10829);
  and g20522 (n10830, n1192, n_10333);
  not g20523 (n_10334, n10830);
  and g20524 (n10831, n1196, n_10334);
  not g20525 (n_10335, n10831);
  and g20526 (n10832, n1200, n_10335);
  not g20527 (n_10336, n10832);
  and g20528 (n10833, n1204, n_10336);
  not g20529 (n_10337, n10833);
  and g20530 (n10834, n1208, n_10337);
  not g20531 (n_10338, n10834);
  and g20532 (n10835, n1212, n_10338);
  not g20533 (n_10339, n10835);
  and g20534 (n10836, n1216, n_10339);
  not g20535 (n_10340, n10836);
  and g20536 (n10837, n1220, n_10340);
  not g20537 (n_10341, n10837);
  and g20538 (n10838, n1224, n_10341);
  not g20539 (n_10342, n10838);
  and g20540 (n10839, n1228, n_10342);
  not g20541 (n_10343, n10839);
  and g20542 (n10840, n1232, n_10343);
  not g20543 (n_10344, n10840);
  and g20544 (n10841, n1236, n_10344);
  not g20545 (n_10345, n10841);
  and g20546 (n10842, n1240, n_10345);
  not g20547 (n_10346, n10842);
  and g20548 (n10843, n1244, n_10346);
  not g20549 (n_10347, n10843);
  and g20550 (n10844, n1248, n_10347);
  not g20551 (n_10348, n10844);
  and g20552 (n10845, n1252, n_10348);
  not g20553 (n_10349, n10845);
  and g20554 (n10846, n1256, n_10349);
  not g20555 (n_10350, n10846);
  and g20556 (n10847, n1260, n_10350);
  not g20557 (n_10351, n10847);
  and g20558 (n10848, n1264, n_10351);
  not g20559 (n_10352, n10848);
  and g20560 (n10849, n1268, n_10352);
  not g20561 (n_10353, n10849);
  and g20562 (n10850, n1272, n_10353);
  not g20563 (n_10354, n10850);
  and g20564 (n10851, n1276, n_10354);
  not g20565 (n_10355, n10851);
  and g20566 (n10852, n1280, n_10355);
  not g20567 (n_10356, n10852);
  and g20568 (n10853, n1284, n_10356);
  not g20569 (n_10357, n10853);
  and g20570 (n10854, n1288, n_10357);
  not g20571 (n_10358, n10854);
  and g20572 (n10855, n1292, n_10358);
  not g20573 (n_10359, n10855);
  and g20574 (n10856, n1296, n_10359);
  not g20575 (n_10360, n10856);
  and g20576 (n10857, n1300, n_10360);
  not g20577 (n_10361, n10857);
  and g20578 (n10858, n1304, n_10361);
  not g20579 (n_10362, n10858);
  and g20580 (n10859, n1308, n_10362);
  not g20581 (n_10363, n10859);
  and g20582 (n10860, n1312, n_10363);
  not g20583 (n_10364, n10860);
  and g20584 (n10861, n1316, n_10364);
  not g20585 (n_10365, n10861);
  and g20586 (n10862, n1320, n_10365);
  not g20587 (n_10366, n10862);
  and g20588 (n10863, n1324, n_10366);
  not g20589 (n_10367, n10863);
  and g20590 (n10864, n1328, n_10367);
  not g20591 (n_10368, n10864);
  and g20592 (n10865, n1332, n_10368);
  not g20593 (n_10369, n10865);
  and g20594 (n10866, n1336, n_10369);
  not g20595 (n_10370, n10866);
  and g20596 (n10867, n1340, n_10370);
  not g20597 (n_10371, n10867);
  and g20598 (n10868, n1344, n_10371);
  not g20599 (n_10372, n10868);
  and g20600 (n10869, n1348, n_10372);
  and g20601 (n10870, \req[112] , n_995);
  not g20602 (n_10373, n10869);
  and g20603 (\grant[112] , n_10373, n10870);
  not g20604 (n_10374, n687);
  and g20605 (n10872, n_10374, n1359);
  not g20606 (n_10375, n10872);
  and g20607 (n10873, n1364, n_10375);
  not g20608 (n_10376, n10873);
  and g20609 (n10874, n1368, n_10376);
  not g20610 (n_10377, n10874);
  and g20611 (n10875, n1372, n_10377);
  not g20612 (n_10378, n10875);
  and g20613 (n10876, n1376, n_10378);
  not g20614 (n_10379, n10876);
  and g20615 (n10877, n1380, n_10379);
  not g20616 (n_10380, n10877);
  and g20617 (n10878, n1384, n_10380);
  not g20618 (n_10381, n10878);
  and g20619 (n10879, n1388, n_10381);
  not g20620 (n_10382, n10879);
  and g20621 (n10880, n1392, n_10382);
  not g20622 (n_10383, n10880);
  and g20623 (n10881, n1396, n_10383);
  not g20624 (n_10384, n10881);
  and g20625 (n10882, n1663, n_10384);
  not g20626 (n_10385, n10882);
  and g20627 (n10883, n392, n_10385);
  not g20628 (n_10386, n10883);
  and g20629 (n10884, n396, n_10386);
  not g20630 (n_10387, n10884);
  and g20631 (n10885, n400, n_10387);
  not g20632 (n_10388, n10885);
  and g20633 (n10886, n404, n_10388);
  not g20634 (n_10389, n10886);
  and g20635 (n10887, n408, n_10389);
  not g20636 (n_10390, n10887);
  and g20637 (n10888, n412, n_10390);
  not g20638 (n_10391, n10888);
  and g20639 (n10889, n416, n_10391);
  not g20640 (n_10392, n10889);
  and g20641 (n10890, n420, n_10392);
  not g20642 (n_10393, n10890);
  and g20643 (n10891, n424, n_10393);
  not g20644 (n_10394, n10891);
  and g20645 (n10892, n428, n_10394);
  not g20646 (n_10395, n10892);
  and g20647 (n10893, n432, n_10395);
  not g20648 (n_10396, n10893);
  and g20649 (n10894, n436, n_10396);
  not g20650 (n_10397, n10894);
  and g20651 (n10895, n440, n_10397);
  not g20652 (n_10398, n10895);
  and g20653 (n10896, n444, n_10398);
  not g20654 (n_10399, n10896);
  and g20655 (n10897, n448, n_10399);
  not g20656 (n_10400, n10897);
  and g20657 (n10898, n452, n_10400);
  not g20658 (n_10401, n10898);
  and g20659 (n10899, n456, n_10401);
  not g20660 (n_10402, n10899);
  and g20661 (n10900, n460, n_10402);
  not g20662 (n_10403, n10900);
  and g20663 (n10901, n464, n_10403);
  not g20664 (n_10404, n10901);
  and g20665 (n10902, n468, n_10404);
  not g20666 (n_10405, n10902);
  and g20667 (n10903, n472, n_10405);
  not g20668 (n_10406, n10903);
  and g20669 (n10904, n476, n_10406);
  not g20670 (n_10407, n10904);
  and g20671 (n10905, n480, n_10407);
  not g20672 (n_10408, n10905);
  and g20673 (n10906, n484, n_10408);
  not g20674 (n_10409, n10906);
  and g20675 (n10907, n488, n_10409);
  not g20676 (n_10410, n10907);
  and g20677 (n10908, n492, n_10410);
  not g20678 (n_10411, n10908);
  and g20679 (n10909, n496, n_10411);
  not g20680 (n_10412, n10909);
  and g20681 (n10910, n500, n_10412);
  not g20682 (n_10413, n10910);
  and g20683 (n10911, n504, n_10413);
  not g20684 (n_10414, n10911);
  and g20685 (n10912, n508, n_10414);
  not g20686 (n_10415, n10912);
  and g20687 (n10913, n512, n_10415);
  not g20688 (n_10416, n10913);
  and g20689 (n10914, n516, n_10416);
  not g20690 (n_10417, n10914);
  and g20691 (n10915, n520, n_10417);
  not g20692 (n_10418, n10915);
  and g20693 (n10916, n524, n_10418);
  not g20694 (n_10419, n10916);
  and g20695 (n10917, n528, n_10419);
  not g20696 (n_10420, n10917);
  and g20697 (n10918, n532, n_10420);
  not g20698 (n_10421, n10918);
  and g20699 (n10919, n536, n_10421);
  not g20700 (n_10422, n10919);
  and g20701 (n10920, n540, n_10422);
  not g20702 (n_10423, n10920);
  and g20703 (n10921, n544, n_10423);
  not g20704 (n_10424, n10921);
  and g20705 (n10922, n548, n_10424);
  not g20706 (n_10425, n10922);
  and g20707 (n10923, n552, n_10425);
  not g20708 (n_10426, n10923);
  and g20709 (n10924, n556, n_10426);
  not g20710 (n_10427, n10924);
  and g20711 (n10925, n560, n_10427);
  not g20712 (n_10428, n10925);
  and g20713 (n10926, n564, n_10428);
  not g20714 (n_10429, n10926);
  and g20715 (n10927, n568, n_10429);
  not g20716 (n_10430, n10927);
  and g20717 (n10928, n572, n_10430);
  not g20718 (n_10431, n10928);
  and g20719 (n10929, n576, n_10431);
  not g20720 (n_10432, n10929);
  and g20721 (n10930, n580, n_10432);
  not g20722 (n_10433, n10930);
  and g20723 (n10931, n584, n_10433);
  not g20724 (n_10434, n10931);
  and g20725 (n10932, n588, n_10434);
  not g20726 (n_10435, n10932);
  and g20727 (n10933, n592, n_10435);
  not g20728 (n_10436, n10933);
  and g20729 (n10934, n596, n_10436);
  not g20730 (n_10437, n10934);
  and g20731 (n10935, n600, n_10437);
  not g20732 (n_10438, n10935);
  and g20733 (n10936, n604, n_10438);
  not g20734 (n_10439, n10936);
  and g20735 (n10937, n608, n_10439);
  not g20736 (n_10440, n10937);
  and g20737 (n10938, n612, n_10440);
  not g20738 (n_10441, n10938);
  and g20739 (n10939, n616, n_10441);
  not g20740 (n_10442, n10939);
  and g20741 (n10940, n620, n_10442);
  not g20742 (n_10443, n10940);
  and g20743 (n10941, n624, n_10443);
  not g20744 (n_10444, n10941);
  and g20745 (n10942, n628, n_10444);
  not g20746 (n_10445, n10942);
  and g20747 (n10943, n632, n_10445);
  not g20748 (n_10446, n10943);
  and g20749 (n10944, n636, n_10446);
  not g20750 (n_10447, n10944);
  and g20751 (n10945, n640, n_10447);
  not g20752 (n_10448, n10945);
  and g20753 (n10946, n644, n_10448);
  not g20754 (n_10449, n10946);
  and g20755 (n10947, n648, n_10449);
  not g20756 (n_10450, n10947);
  and g20757 (n10948, n652, n_10450);
  not g20758 (n_10451, n10948);
  and g20759 (n10949, n656, n_10451);
  not g20760 (n_10452, n10949);
  and g20761 (n10950, n660, n_10452);
  not g20762 (n_10453, n10950);
  and g20763 (n10951, n664, n_10453);
  not g20764 (n_10454, n10951);
  and g20765 (n10952, n668, n_10454);
  not g20766 (n_10455, n10952);
  and g20767 (n10953, n672, n_10455);
  not g20768 (n_10456, n10953);
  and g20769 (n10954, n676, n_10456);
  not g20770 (n_10457, n10954);
  and g20771 (n10955, n680, n_10457);
  and g20772 (n10956, \req[113] , n_528);
  not g20773 (n_10458, n10955);
  and g20774 (\grant[113] , n_10458, n10956);
  not g20775 (n_10459, n1026);
  and g20776 (n10958, n691, n_10459);
  not g20777 (n_10460, n10958);
  and g20778 (n10959, n696, n_10460);
  not g20779 (n_10461, n10959);
  and g20780 (n10960, n700, n_10461);
  not g20781 (n_10462, n10960);
  and g20782 (n10961, n704, n_10462);
  not g20783 (n_10463, n10961);
  and g20784 (n10962, n708, n_10463);
  not g20785 (n_10464, n10962);
  and g20786 (n10963, n712, n_10464);
  not g20787 (n_10465, n10963);
  and g20788 (n10964, n716, n_10465);
  not g20789 (n_10466, n10964);
  and g20790 (n10965, n720, n_10466);
  not g20791 (n_10467, n10965);
  and g20792 (n10966, n1484, n_10467);
  not g20793 (n_10468, n10966);
  and g20794 (n10967, n1486, n_10468);
  not g20795 (n_10469, n10967);
  and g20796 (n10968, n1750, n_10469);
  not g20797 (n_10470, n10968);
  and g20798 (n10969, n731, n_10470);
  not g20799 (n_10471, n10969);
  and g20800 (n10970, n735, n_10471);
  not g20801 (n_10472, n10970);
  and g20802 (n10971, n739, n_10472);
  not g20803 (n_10473, n10971);
  and g20804 (n10972, n743, n_10473);
  not g20805 (n_10474, n10972);
  and g20806 (n10973, n747, n_10474);
  not g20807 (n_10475, n10973);
  and g20808 (n10974, n751, n_10475);
  not g20809 (n_10476, n10974);
  and g20810 (n10975, n755, n_10476);
  not g20811 (n_10477, n10975);
  and g20812 (n10976, n759, n_10477);
  not g20813 (n_10478, n10976);
  and g20814 (n10977, n763, n_10478);
  not g20815 (n_10479, n10977);
  and g20816 (n10978, n767, n_10479);
  not g20817 (n_10480, n10978);
  and g20818 (n10979, n771, n_10480);
  not g20819 (n_10481, n10979);
  and g20820 (n10980, n775, n_10481);
  not g20821 (n_10482, n10980);
  and g20822 (n10981, n779, n_10482);
  not g20823 (n_10483, n10981);
  and g20824 (n10982, n783, n_10483);
  not g20825 (n_10484, n10982);
  and g20826 (n10983, n787, n_10484);
  not g20827 (n_10485, n10983);
  and g20828 (n10984, n791, n_10485);
  not g20829 (n_10486, n10984);
  and g20830 (n10985, n795, n_10486);
  not g20831 (n_10487, n10985);
  and g20832 (n10986, n799, n_10487);
  not g20833 (n_10488, n10986);
  and g20834 (n10987, n803, n_10488);
  not g20835 (n_10489, n10987);
  and g20836 (n10988, n807, n_10489);
  not g20837 (n_10490, n10988);
  and g20838 (n10989, n811, n_10490);
  not g20839 (n_10491, n10989);
  and g20840 (n10990, n815, n_10491);
  not g20841 (n_10492, n10990);
  and g20842 (n10991, n819, n_10492);
  not g20843 (n_10493, n10991);
  and g20844 (n10992, n823, n_10493);
  not g20845 (n_10494, n10992);
  and g20846 (n10993, n827, n_10494);
  not g20847 (n_10495, n10993);
  and g20848 (n10994, n831, n_10495);
  not g20849 (n_10496, n10994);
  and g20850 (n10995, n835, n_10496);
  not g20851 (n_10497, n10995);
  and g20852 (n10996, n839, n_10497);
  not g20853 (n_10498, n10996);
  and g20854 (n10997, n843, n_10498);
  not g20855 (n_10499, n10997);
  and g20856 (n10998, n847, n_10499);
  not g20857 (n_10500, n10998);
  and g20858 (n10999, n851, n_10500);
  not g20859 (n_10501, n10999);
  and g20860 (n11000, n855, n_10501);
  not g20861 (n_10502, n11000);
  and g20862 (n11001, n859, n_10502);
  not g20863 (n_10503, n11001);
  and g20864 (n11002, n863, n_10503);
  not g20865 (n_10504, n11002);
  and g20866 (n11003, n867, n_10504);
  not g20867 (n_10505, n11003);
  and g20868 (n11004, n871, n_10505);
  not g20869 (n_10506, n11004);
  and g20870 (n11005, n875, n_10506);
  not g20871 (n_10507, n11005);
  and g20872 (n11006, n879, n_10507);
  not g20873 (n_10508, n11006);
  and g20874 (n11007, n883, n_10508);
  not g20875 (n_10509, n11007);
  and g20876 (n11008, n887, n_10509);
  not g20877 (n_10510, n11008);
  and g20878 (n11009, n891, n_10510);
  not g20879 (n_10511, n11009);
  and g20880 (n11010, n895, n_10511);
  not g20881 (n_10512, n11010);
  and g20882 (n11011, n899, n_10512);
  not g20883 (n_10513, n11011);
  and g20884 (n11012, n903, n_10513);
  not g20885 (n_10514, n11012);
  and g20886 (n11013, n907, n_10514);
  not g20887 (n_10515, n11013);
  and g20888 (n11014, n911, n_10515);
  not g20889 (n_10516, n11014);
  and g20890 (n11015, n915, n_10516);
  not g20891 (n_10517, n11015);
  and g20892 (n11016, n919, n_10517);
  not g20893 (n_10518, n11016);
  and g20894 (n11017, n923, n_10518);
  not g20895 (n_10519, n11017);
  and g20896 (n11018, n927, n_10519);
  not g20897 (n_10520, n11018);
  and g20898 (n11019, n931, n_10520);
  not g20899 (n_10521, n11019);
  and g20900 (n11020, n935, n_10521);
  not g20901 (n_10522, n11020);
  and g20902 (n11021, n939, n_10522);
  not g20903 (n_10523, n11021);
  and g20904 (n11022, n943, n_10523);
  not g20905 (n_10524, n11022);
  and g20906 (n11023, n947, n_10524);
  not g20907 (n_10525, n11023);
  and g20908 (n11024, n951, n_10525);
  not g20909 (n_10526, n11024);
  and g20910 (n11025, n955, n_10526);
  not g20911 (n_10527, n11025);
  and g20912 (n11026, n959, n_10527);
  not g20913 (n_10528, n11026);
  and g20914 (n11027, n963, n_10528);
  not g20915 (n_10529, n11027);
  and g20916 (n11028, n967, n_10529);
  not g20917 (n_10530, n11028);
  and g20918 (n11029, n971, n_10530);
  not g20919 (n_10531, n11029);
  and g20920 (n11030, n975, n_10531);
  not g20921 (n_10532, n11030);
  and g20922 (n11031, n979, n_10532);
  not g20923 (n_10533, n11031);
  and g20924 (n11032, n983, n_10533);
  not g20925 (n_10534, n11032);
  and g20926 (n11033, n987, n_10534);
  not g20927 (n_10535, n11033);
  and g20928 (n11034, n991, n_10535);
  not g20929 (n_10536, n11034);
  and g20930 (n11035, n995, n_10536);
  not g20931 (n_10537, n11035);
  and g20932 (n11036, n999, n_10537);
  not g20933 (n_10538, n11036);
  and g20934 (n11037, n1003, n_10538);
  not g20935 (n_10539, n11037);
  and g20936 (n11038, n1007, n_10539);
  not g20937 (n_10540, n11038);
  and g20938 (n11039, n1011, n_10540);
  not g20939 (n_10541, n11039);
  and g20940 (n11040, n1015, n_10541);
  not g20941 (n_10542, n11040);
  and g20942 (n11041, n1019, n_10542);
  and g20943 (n11042, \req[114] , n_821);
  not g20944 (n_10543, n11041);
  and g20945 (\grant[114] , n_10543, n11042);
  not g20946 (n_10544, n1363);
  and g20947 (n11044, n1030, n_10544);
  not g20948 (n_10545, n11044);
  and g20949 (n11045, n1035, n_10545);
  not g20950 (n_10546, n11045);
  and g20951 (n11046, n1039, n_10546);
  not g20952 (n_10547, n11046);
  and g20953 (n11047, n1043, n_10547);
  not g20954 (n_10548, n11047);
  and g20955 (n11048, n1047, n_10548);
  not g20956 (n_10549, n11048);
  and g20957 (n11049, n1051, n_10549);
  not g20958 (n_10550, n11049);
  and g20959 (n11050, n1055, n_10550);
  not g20960 (n_10551, n11050);
  and g20961 (n11051, n1059, n_10551);
  not g20962 (n_10552, n11051);
  and g20963 (n11052, n1574, n_10552);
  not g20964 (n_10553, n11052);
  and g20965 (n11053, n1576, n_10553);
  not g20966 (n_10554, n11053);
  and g20967 (n11054, n1837, n_10554);
  not g20968 (n_10555, n11054);
  and g20969 (n11055, n1068, n_10555);
  not g20970 (n_10556, n11055);
  and g20971 (n11056, n1072, n_10556);
  not g20972 (n_10557, n11056);
  and g20973 (n11057, n1076, n_10557);
  not g20974 (n_10558, n11057);
  and g20975 (n11058, n1080, n_10558);
  not g20976 (n_10559, n11058);
  and g20977 (n11059, n1084, n_10559);
  not g20978 (n_10560, n11059);
  and g20979 (n11060, n1088, n_10560);
  not g20980 (n_10561, n11060);
  and g20981 (n11061, n1092, n_10561);
  not g20982 (n_10562, n11061);
  and g20983 (n11062, n1096, n_10562);
  not g20984 (n_10563, n11062);
  and g20985 (n11063, n1100, n_10563);
  not g20986 (n_10564, n11063);
  and g20987 (n11064, n1104, n_10564);
  not g20988 (n_10565, n11064);
  and g20989 (n11065, n1108, n_10565);
  not g20990 (n_10566, n11065);
  and g20991 (n11066, n1112, n_10566);
  not g20992 (n_10567, n11066);
  and g20993 (n11067, n1116, n_10567);
  not g20994 (n_10568, n11067);
  and g20995 (n11068, n1120, n_10568);
  not g20996 (n_10569, n11068);
  and g20997 (n11069, n1124, n_10569);
  not g20998 (n_10570, n11069);
  and g20999 (n11070, n1128, n_10570);
  not g21000 (n_10571, n11070);
  and g21001 (n11071, n1132, n_10571);
  not g21002 (n_10572, n11071);
  and g21003 (n11072, n1136, n_10572);
  not g21004 (n_10573, n11072);
  and g21005 (n11073, n1140, n_10573);
  not g21006 (n_10574, n11073);
  and g21007 (n11074, n1144, n_10574);
  not g21008 (n_10575, n11074);
  and g21009 (n11075, n1148, n_10575);
  not g21010 (n_10576, n11075);
  and g21011 (n11076, n1152, n_10576);
  not g21012 (n_10577, n11076);
  and g21013 (n11077, n1156, n_10577);
  not g21014 (n_10578, n11077);
  and g21015 (n11078, n1160, n_10578);
  not g21016 (n_10579, n11078);
  and g21017 (n11079, n1164, n_10579);
  not g21018 (n_10580, n11079);
  and g21019 (n11080, n1168, n_10580);
  not g21020 (n_10581, n11080);
  and g21021 (n11081, n1172, n_10581);
  not g21022 (n_10582, n11081);
  and g21023 (n11082, n1176, n_10582);
  not g21024 (n_10583, n11082);
  and g21025 (n11083, n1180, n_10583);
  not g21026 (n_10584, n11083);
  and g21027 (n11084, n1184, n_10584);
  not g21028 (n_10585, n11084);
  and g21029 (n11085, n1188, n_10585);
  not g21030 (n_10586, n11085);
  and g21031 (n11086, n1192, n_10586);
  not g21032 (n_10587, n11086);
  and g21033 (n11087, n1196, n_10587);
  not g21034 (n_10588, n11087);
  and g21035 (n11088, n1200, n_10588);
  not g21036 (n_10589, n11088);
  and g21037 (n11089, n1204, n_10589);
  not g21038 (n_10590, n11089);
  and g21039 (n11090, n1208, n_10590);
  not g21040 (n_10591, n11090);
  and g21041 (n11091, n1212, n_10591);
  not g21042 (n_10592, n11091);
  and g21043 (n11092, n1216, n_10592);
  not g21044 (n_10593, n11092);
  and g21045 (n11093, n1220, n_10593);
  not g21046 (n_10594, n11093);
  and g21047 (n11094, n1224, n_10594);
  not g21048 (n_10595, n11094);
  and g21049 (n11095, n1228, n_10595);
  not g21050 (n_10596, n11095);
  and g21051 (n11096, n1232, n_10596);
  not g21052 (n_10597, n11096);
  and g21053 (n11097, n1236, n_10597);
  not g21054 (n_10598, n11097);
  and g21055 (n11098, n1240, n_10598);
  not g21056 (n_10599, n11098);
  and g21057 (n11099, n1244, n_10599);
  not g21058 (n_10600, n11099);
  and g21059 (n11100, n1248, n_10600);
  not g21060 (n_10601, n11100);
  and g21061 (n11101, n1252, n_10601);
  not g21062 (n_10602, n11101);
  and g21063 (n11102, n1256, n_10602);
  not g21064 (n_10603, n11102);
  and g21065 (n11103, n1260, n_10603);
  not g21066 (n_10604, n11103);
  and g21067 (n11104, n1264, n_10604);
  not g21068 (n_10605, n11104);
  and g21069 (n11105, n1268, n_10605);
  not g21070 (n_10606, n11105);
  and g21071 (n11106, n1272, n_10606);
  not g21072 (n_10607, n11106);
  and g21073 (n11107, n1276, n_10607);
  not g21074 (n_10608, n11107);
  and g21075 (n11108, n1280, n_10608);
  not g21076 (n_10609, n11108);
  and g21077 (n11109, n1284, n_10609);
  not g21078 (n_10610, n11109);
  and g21079 (n11110, n1288, n_10610);
  not g21080 (n_10611, n11110);
  and g21081 (n11111, n1292, n_10611);
  not g21082 (n_10612, n11111);
  and g21083 (n11112, n1296, n_10612);
  not g21084 (n_10613, n11112);
  and g21085 (n11113, n1300, n_10613);
  not g21086 (n_10614, n11113);
  and g21087 (n11114, n1304, n_10614);
  not g21088 (n_10615, n11114);
  and g21089 (n11115, n1308, n_10615);
  not g21090 (n_10616, n11115);
  and g21091 (n11116, n1312, n_10616);
  not g21092 (n_10617, n11116);
  and g21093 (n11117, n1316, n_10617);
  not g21094 (n_10618, n11117);
  and g21095 (n11118, n1320, n_10618);
  not g21096 (n_10619, n11118);
  and g21097 (n11119, n1324, n_10619);
  not g21098 (n_10620, n11119);
  and g21099 (n11120, n1328, n_10620);
  not g21100 (n_10621, n11120);
  and g21101 (n11121, n1332, n_10621);
  not g21102 (n_10622, n11121);
  and g21103 (n11122, n1336, n_10622);
  not g21104 (n_10623, n11122);
  and g21105 (n11123, n1340, n_10623);
  not g21106 (n_10624, n11123);
  and g21107 (n11124, n1344, n_10624);
  not g21108 (n_10625, n11124);
  and g21109 (n11125, n1348, n_10625);
  not g21110 (n_10626, n11125);
  and g21111 (n11126, n1352, n_10626);
  not g21112 (n_10627, n11126);
  and g21113 (n11127, n1356, n_10627);
  and g21114 (n11128, \req[115] , n_999);
  not g21115 (n_10628, n11127);
  and g21116 (\grant[115] , n_10628, n11128);
  not g21117 (n_10629, n695);
  and g21118 (n11130, n_10629, n1367);
  not g21119 (n_10630, n11130);
  and g21120 (n11131, n1372, n_10630);
  not g21121 (n_10631, n11131);
  and g21122 (n11132, n1376, n_10631);
  not g21123 (n_10632, n11132);
  and g21124 (n11133, n1380, n_10632);
  not g21125 (n_10633, n11133);
  and g21126 (n11134, n1384, n_10633);
  not g21127 (n_10634, n11134);
  and g21128 (n11135, n1388, n_10634);
  not g21129 (n_10635, n11135);
  and g21130 (n11136, n1392, n_10635);
  not g21131 (n_10636, n11136);
  and g21132 (n11137, n1396, n_10636);
  not g21133 (n_10637, n11137);
  and g21134 (n11138, n1663, n_10637);
  not g21135 (n_10638, n11138);
  and g21136 (n11139, n392, n_10638);
  not g21137 (n_10639, n11139);
  and g21138 (n11140, n396, n_10639);
  not g21139 (n_10640, n11140);
  and g21140 (n11141, n400, n_10640);
  not g21141 (n_10641, n11141);
  and g21142 (n11142, n404, n_10641);
  not g21143 (n_10642, n11142);
  and g21144 (n11143, n408, n_10642);
  not g21145 (n_10643, n11143);
  and g21146 (n11144, n412, n_10643);
  not g21147 (n_10644, n11144);
  and g21148 (n11145, n416, n_10644);
  not g21149 (n_10645, n11145);
  and g21150 (n11146, n420, n_10645);
  not g21151 (n_10646, n11146);
  and g21152 (n11147, n424, n_10646);
  not g21153 (n_10647, n11147);
  and g21154 (n11148, n428, n_10647);
  not g21155 (n_10648, n11148);
  and g21156 (n11149, n432, n_10648);
  not g21157 (n_10649, n11149);
  and g21158 (n11150, n436, n_10649);
  not g21159 (n_10650, n11150);
  and g21160 (n11151, n440, n_10650);
  not g21161 (n_10651, n11151);
  and g21162 (n11152, n444, n_10651);
  not g21163 (n_10652, n11152);
  and g21164 (n11153, n448, n_10652);
  not g21165 (n_10653, n11153);
  and g21166 (n11154, n452, n_10653);
  not g21167 (n_10654, n11154);
  and g21168 (n11155, n456, n_10654);
  not g21169 (n_10655, n11155);
  and g21170 (n11156, n460, n_10655);
  not g21171 (n_10656, n11156);
  and g21172 (n11157, n464, n_10656);
  not g21173 (n_10657, n11157);
  and g21174 (n11158, n468, n_10657);
  not g21175 (n_10658, n11158);
  and g21176 (n11159, n472, n_10658);
  not g21177 (n_10659, n11159);
  and g21178 (n11160, n476, n_10659);
  not g21179 (n_10660, n11160);
  and g21180 (n11161, n480, n_10660);
  not g21181 (n_10661, n11161);
  and g21182 (n11162, n484, n_10661);
  not g21183 (n_10662, n11162);
  and g21184 (n11163, n488, n_10662);
  not g21185 (n_10663, n11163);
  and g21186 (n11164, n492, n_10663);
  not g21187 (n_10664, n11164);
  and g21188 (n11165, n496, n_10664);
  not g21189 (n_10665, n11165);
  and g21190 (n11166, n500, n_10665);
  not g21191 (n_10666, n11166);
  and g21192 (n11167, n504, n_10666);
  not g21193 (n_10667, n11167);
  and g21194 (n11168, n508, n_10667);
  not g21195 (n_10668, n11168);
  and g21196 (n11169, n512, n_10668);
  not g21197 (n_10669, n11169);
  and g21198 (n11170, n516, n_10669);
  not g21199 (n_10670, n11170);
  and g21200 (n11171, n520, n_10670);
  not g21201 (n_10671, n11171);
  and g21202 (n11172, n524, n_10671);
  not g21203 (n_10672, n11172);
  and g21204 (n11173, n528, n_10672);
  not g21205 (n_10673, n11173);
  and g21206 (n11174, n532, n_10673);
  not g21207 (n_10674, n11174);
  and g21208 (n11175, n536, n_10674);
  not g21209 (n_10675, n11175);
  and g21210 (n11176, n540, n_10675);
  not g21211 (n_10676, n11176);
  and g21212 (n11177, n544, n_10676);
  not g21213 (n_10677, n11177);
  and g21214 (n11178, n548, n_10677);
  not g21215 (n_10678, n11178);
  and g21216 (n11179, n552, n_10678);
  not g21217 (n_10679, n11179);
  and g21218 (n11180, n556, n_10679);
  not g21219 (n_10680, n11180);
  and g21220 (n11181, n560, n_10680);
  not g21221 (n_10681, n11181);
  and g21222 (n11182, n564, n_10681);
  not g21223 (n_10682, n11182);
  and g21224 (n11183, n568, n_10682);
  not g21225 (n_10683, n11183);
  and g21226 (n11184, n572, n_10683);
  not g21227 (n_10684, n11184);
  and g21228 (n11185, n576, n_10684);
  not g21229 (n_10685, n11185);
  and g21230 (n11186, n580, n_10685);
  not g21231 (n_10686, n11186);
  and g21232 (n11187, n584, n_10686);
  not g21233 (n_10687, n11187);
  and g21234 (n11188, n588, n_10687);
  not g21235 (n_10688, n11188);
  and g21236 (n11189, n592, n_10688);
  not g21237 (n_10689, n11189);
  and g21238 (n11190, n596, n_10689);
  not g21239 (n_10690, n11190);
  and g21240 (n11191, n600, n_10690);
  not g21241 (n_10691, n11191);
  and g21242 (n11192, n604, n_10691);
  not g21243 (n_10692, n11192);
  and g21244 (n11193, n608, n_10692);
  not g21245 (n_10693, n11193);
  and g21246 (n11194, n612, n_10693);
  not g21247 (n_10694, n11194);
  and g21248 (n11195, n616, n_10694);
  not g21249 (n_10695, n11195);
  and g21250 (n11196, n620, n_10695);
  not g21251 (n_10696, n11196);
  and g21252 (n11197, n624, n_10696);
  not g21253 (n_10697, n11197);
  and g21254 (n11198, n628, n_10697);
  not g21255 (n_10698, n11198);
  and g21256 (n11199, n632, n_10698);
  not g21257 (n_10699, n11199);
  and g21258 (n11200, n636, n_10699);
  not g21259 (n_10700, n11200);
  and g21260 (n11201, n640, n_10700);
  not g21261 (n_10701, n11201);
  and g21262 (n11202, n644, n_10701);
  not g21263 (n_10702, n11202);
  and g21264 (n11203, n648, n_10702);
  not g21265 (n_10703, n11203);
  and g21266 (n11204, n652, n_10703);
  not g21267 (n_10704, n11204);
  and g21268 (n11205, n656, n_10704);
  not g21269 (n_10705, n11205);
  and g21270 (n11206, n660, n_10705);
  not g21271 (n_10706, n11206);
  and g21272 (n11207, n664, n_10706);
  not g21273 (n_10707, n11207);
  and g21274 (n11208, n668, n_10707);
  not g21275 (n_10708, n11208);
  and g21276 (n11209, n672, n_10708);
  not g21277 (n_10709, n11209);
  and g21278 (n11210, n676, n_10709);
  not g21279 (n_10710, n11210);
  and g21280 (n11211, n680, n_10710);
  not g21281 (n_10711, n11211);
  and g21282 (n11212, n684, n_10711);
  not g21283 (n_10712, n11212);
  and g21284 (n11213, n688, n_10712);
  and g21285 (n11214, \req[116] , n_542);
  not g21286 (n_10713, n11213);
  and g21287 (\grant[116] , n_10713, n11214);
  not g21288 (n_10714, n1034);
  and g21289 (n11216, n699, n_10714);
  not g21290 (n_10715, n11216);
  and g21291 (n11217, n704, n_10715);
  not g21292 (n_10716, n11217);
  and g21293 (n11218, n708, n_10716);
  not g21294 (n_10717, n11218);
  and g21295 (n11219, n712, n_10717);
  not g21296 (n_10718, n11219);
  and g21297 (n11220, n716, n_10718);
  not g21298 (n_10719, n11220);
  and g21299 (n11221, n720, n_10719);
  not g21300 (n_10720, n11221);
  and g21301 (n11222, n1484, n_10720);
  not g21302 (n_10721, n11222);
  and g21303 (n11223, n1486, n_10721);
  not g21304 (n_10722, n11223);
  and g21305 (n11224, n1750, n_10722);
  not g21306 (n_10723, n11224);
  and g21307 (n11225, n731, n_10723);
  not g21308 (n_10724, n11225);
  and g21309 (n11226, n735, n_10724);
  not g21310 (n_10725, n11226);
  and g21311 (n11227, n739, n_10725);
  not g21312 (n_10726, n11227);
  and g21313 (n11228, n743, n_10726);
  not g21314 (n_10727, n11228);
  and g21315 (n11229, n747, n_10727);
  not g21316 (n_10728, n11229);
  and g21317 (n11230, n751, n_10728);
  not g21318 (n_10729, n11230);
  and g21319 (n11231, n755, n_10729);
  not g21320 (n_10730, n11231);
  and g21321 (n11232, n759, n_10730);
  not g21322 (n_10731, n11232);
  and g21323 (n11233, n763, n_10731);
  not g21324 (n_10732, n11233);
  and g21325 (n11234, n767, n_10732);
  not g21326 (n_10733, n11234);
  and g21327 (n11235, n771, n_10733);
  not g21328 (n_10734, n11235);
  and g21329 (n11236, n775, n_10734);
  not g21330 (n_10735, n11236);
  and g21331 (n11237, n779, n_10735);
  not g21332 (n_10736, n11237);
  and g21333 (n11238, n783, n_10736);
  not g21334 (n_10737, n11238);
  and g21335 (n11239, n787, n_10737);
  not g21336 (n_10738, n11239);
  and g21337 (n11240, n791, n_10738);
  not g21338 (n_10739, n11240);
  and g21339 (n11241, n795, n_10739);
  not g21340 (n_10740, n11241);
  and g21341 (n11242, n799, n_10740);
  not g21342 (n_10741, n11242);
  and g21343 (n11243, n803, n_10741);
  not g21344 (n_10742, n11243);
  and g21345 (n11244, n807, n_10742);
  not g21346 (n_10743, n11244);
  and g21347 (n11245, n811, n_10743);
  not g21348 (n_10744, n11245);
  and g21349 (n11246, n815, n_10744);
  not g21350 (n_10745, n11246);
  and g21351 (n11247, n819, n_10745);
  not g21352 (n_10746, n11247);
  and g21353 (n11248, n823, n_10746);
  not g21354 (n_10747, n11248);
  and g21355 (n11249, n827, n_10747);
  not g21356 (n_10748, n11249);
  and g21357 (n11250, n831, n_10748);
  not g21358 (n_10749, n11250);
  and g21359 (n11251, n835, n_10749);
  not g21360 (n_10750, n11251);
  and g21361 (n11252, n839, n_10750);
  not g21362 (n_10751, n11252);
  and g21363 (n11253, n843, n_10751);
  not g21364 (n_10752, n11253);
  and g21365 (n11254, n847, n_10752);
  not g21366 (n_10753, n11254);
  and g21367 (n11255, n851, n_10753);
  not g21368 (n_10754, n11255);
  and g21369 (n11256, n855, n_10754);
  not g21370 (n_10755, n11256);
  and g21371 (n11257, n859, n_10755);
  not g21372 (n_10756, n11257);
  and g21373 (n11258, n863, n_10756);
  not g21374 (n_10757, n11258);
  and g21375 (n11259, n867, n_10757);
  not g21376 (n_10758, n11259);
  and g21377 (n11260, n871, n_10758);
  not g21378 (n_10759, n11260);
  and g21379 (n11261, n875, n_10759);
  not g21380 (n_10760, n11261);
  and g21381 (n11262, n879, n_10760);
  not g21382 (n_10761, n11262);
  and g21383 (n11263, n883, n_10761);
  not g21384 (n_10762, n11263);
  and g21385 (n11264, n887, n_10762);
  not g21386 (n_10763, n11264);
  and g21387 (n11265, n891, n_10763);
  not g21388 (n_10764, n11265);
  and g21389 (n11266, n895, n_10764);
  not g21390 (n_10765, n11266);
  and g21391 (n11267, n899, n_10765);
  not g21392 (n_10766, n11267);
  and g21393 (n11268, n903, n_10766);
  not g21394 (n_10767, n11268);
  and g21395 (n11269, n907, n_10767);
  not g21396 (n_10768, n11269);
  and g21397 (n11270, n911, n_10768);
  not g21398 (n_10769, n11270);
  and g21399 (n11271, n915, n_10769);
  not g21400 (n_10770, n11271);
  and g21401 (n11272, n919, n_10770);
  not g21402 (n_10771, n11272);
  and g21403 (n11273, n923, n_10771);
  not g21404 (n_10772, n11273);
  and g21405 (n11274, n927, n_10772);
  not g21406 (n_10773, n11274);
  and g21407 (n11275, n931, n_10773);
  not g21408 (n_10774, n11275);
  and g21409 (n11276, n935, n_10774);
  not g21410 (n_10775, n11276);
  and g21411 (n11277, n939, n_10775);
  not g21412 (n_10776, n11277);
  and g21413 (n11278, n943, n_10776);
  not g21414 (n_10777, n11278);
  and g21415 (n11279, n947, n_10777);
  not g21416 (n_10778, n11279);
  and g21417 (n11280, n951, n_10778);
  not g21418 (n_10779, n11280);
  and g21419 (n11281, n955, n_10779);
  not g21420 (n_10780, n11281);
  and g21421 (n11282, n959, n_10780);
  not g21422 (n_10781, n11282);
  and g21423 (n11283, n963, n_10781);
  not g21424 (n_10782, n11283);
  and g21425 (n11284, n967, n_10782);
  not g21426 (n_10783, n11284);
  and g21427 (n11285, n971, n_10783);
  not g21428 (n_10784, n11285);
  and g21429 (n11286, n975, n_10784);
  not g21430 (n_10785, n11286);
  and g21431 (n11287, n979, n_10785);
  not g21432 (n_10786, n11287);
  and g21433 (n11288, n983, n_10786);
  not g21434 (n_10787, n11288);
  and g21435 (n11289, n987, n_10787);
  not g21436 (n_10788, n11289);
  and g21437 (n11290, n991, n_10788);
  not g21438 (n_10789, n11290);
  and g21439 (n11291, n995, n_10789);
  not g21440 (n_10790, n11291);
  and g21441 (n11292, n999, n_10790);
  not g21442 (n_10791, n11292);
  and g21443 (n11293, n1003, n_10791);
  not g21444 (n_10792, n11293);
  and g21445 (n11294, n1007, n_10792);
  not g21446 (n_10793, n11294);
  and g21447 (n11295, n1011, n_10793);
  not g21448 (n_10794, n11295);
  and g21449 (n11296, n1015, n_10794);
  not g21450 (n_10795, n11296);
  and g21451 (n11297, n1019, n_10795);
  not g21452 (n_10796, n11297);
  and g21453 (n11298, n1023, n_10796);
  not g21454 (n_10797, n11298);
  and g21455 (n11299, n1027, n_10797);
  and g21456 (n11300, \req[117] , n_827);
  not g21457 (n_10798, n11299);
  and g21458 (\grant[117] , n_10798, n11300);
  not g21459 (n_10799, n1371);
  and g21460 (n11302, n1038, n_10799);
  not g21461 (n_10800, n11302);
  and g21462 (n11303, n1043, n_10800);
  not g21463 (n_10801, n11303);
  and g21464 (n11304, n1047, n_10801);
  not g21465 (n_10802, n11304);
  and g21466 (n11305, n1051, n_10802);
  not g21467 (n_10803, n11305);
  and g21468 (n11306, n1055, n_10803);
  not g21469 (n_10804, n11306);
  and g21470 (n11307, n1059, n_10804);
  not g21471 (n_10805, n11307);
  and g21472 (n11308, n1574, n_10805);
  not g21473 (n_10806, n11308);
  and g21474 (n11309, n1576, n_10806);
  not g21475 (n_10807, n11309);
  and g21476 (n11310, n1837, n_10807);
  not g21477 (n_10808, n11310);
  and g21478 (n11311, n1068, n_10808);
  not g21479 (n_10809, n11311);
  and g21480 (n11312, n1072, n_10809);
  not g21481 (n_10810, n11312);
  and g21482 (n11313, n1076, n_10810);
  not g21483 (n_10811, n11313);
  and g21484 (n11314, n1080, n_10811);
  not g21485 (n_10812, n11314);
  and g21486 (n11315, n1084, n_10812);
  not g21487 (n_10813, n11315);
  and g21488 (n11316, n1088, n_10813);
  not g21489 (n_10814, n11316);
  and g21490 (n11317, n1092, n_10814);
  not g21491 (n_10815, n11317);
  and g21492 (n11318, n1096, n_10815);
  not g21493 (n_10816, n11318);
  and g21494 (n11319, n1100, n_10816);
  not g21495 (n_10817, n11319);
  and g21496 (n11320, n1104, n_10817);
  not g21497 (n_10818, n11320);
  and g21498 (n11321, n1108, n_10818);
  not g21499 (n_10819, n11321);
  and g21500 (n11322, n1112, n_10819);
  not g21501 (n_10820, n11322);
  and g21502 (n11323, n1116, n_10820);
  not g21503 (n_10821, n11323);
  and g21504 (n11324, n1120, n_10821);
  not g21505 (n_10822, n11324);
  and g21506 (n11325, n1124, n_10822);
  not g21507 (n_10823, n11325);
  and g21508 (n11326, n1128, n_10823);
  not g21509 (n_10824, n11326);
  and g21510 (n11327, n1132, n_10824);
  not g21511 (n_10825, n11327);
  and g21512 (n11328, n1136, n_10825);
  not g21513 (n_10826, n11328);
  and g21514 (n11329, n1140, n_10826);
  not g21515 (n_10827, n11329);
  and g21516 (n11330, n1144, n_10827);
  not g21517 (n_10828, n11330);
  and g21518 (n11331, n1148, n_10828);
  not g21519 (n_10829, n11331);
  and g21520 (n11332, n1152, n_10829);
  not g21521 (n_10830, n11332);
  and g21522 (n11333, n1156, n_10830);
  not g21523 (n_10831, n11333);
  and g21524 (n11334, n1160, n_10831);
  not g21525 (n_10832, n11334);
  and g21526 (n11335, n1164, n_10832);
  not g21527 (n_10833, n11335);
  and g21528 (n11336, n1168, n_10833);
  not g21529 (n_10834, n11336);
  and g21530 (n11337, n1172, n_10834);
  not g21531 (n_10835, n11337);
  and g21532 (n11338, n1176, n_10835);
  not g21533 (n_10836, n11338);
  and g21534 (n11339, n1180, n_10836);
  not g21535 (n_10837, n11339);
  and g21536 (n11340, n1184, n_10837);
  not g21537 (n_10838, n11340);
  and g21538 (n11341, n1188, n_10838);
  not g21539 (n_10839, n11341);
  and g21540 (n11342, n1192, n_10839);
  not g21541 (n_10840, n11342);
  and g21542 (n11343, n1196, n_10840);
  not g21543 (n_10841, n11343);
  and g21544 (n11344, n1200, n_10841);
  not g21545 (n_10842, n11344);
  and g21546 (n11345, n1204, n_10842);
  not g21547 (n_10843, n11345);
  and g21548 (n11346, n1208, n_10843);
  not g21549 (n_10844, n11346);
  and g21550 (n11347, n1212, n_10844);
  not g21551 (n_10845, n11347);
  and g21552 (n11348, n1216, n_10845);
  not g21553 (n_10846, n11348);
  and g21554 (n11349, n1220, n_10846);
  not g21555 (n_10847, n11349);
  and g21556 (n11350, n1224, n_10847);
  not g21557 (n_10848, n11350);
  and g21558 (n11351, n1228, n_10848);
  not g21559 (n_10849, n11351);
  and g21560 (n11352, n1232, n_10849);
  not g21561 (n_10850, n11352);
  and g21562 (n11353, n1236, n_10850);
  not g21563 (n_10851, n11353);
  and g21564 (n11354, n1240, n_10851);
  not g21565 (n_10852, n11354);
  and g21566 (n11355, n1244, n_10852);
  not g21567 (n_10853, n11355);
  and g21568 (n11356, n1248, n_10853);
  not g21569 (n_10854, n11356);
  and g21570 (n11357, n1252, n_10854);
  not g21571 (n_10855, n11357);
  and g21572 (n11358, n1256, n_10855);
  not g21573 (n_10856, n11358);
  and g21574 (n11359, n1260, n_10856);
  not g21575 (n_10857, n11359);
  and g21576 (n11360, n1264, n_10857);
  not g21577 (n_10858, n11360);
  and g21578 (n11361, n1268, n_10858);
  not g21579 (n_10859, n11361);
  and g21580 (n11362, n1272, n_10859);
  not g21581 (n_10860, n11362);
  and g21582 (n11363, n1276, n_10860);
  not g21583 (n_10861, n11363);
  and g21584 (n11364, n1280, n_10861);
  not g21585 (n_10862, n11364);
  and g21586 (n11365, n1284, n_10862);
  not g21587 (n_10863, n11365);
  and g21588 (n11366, n1288, n_10863);
  not g21589 (n_10864, n11366);
  and g21590 (n11367, n1292, n_10864);
  not g21591 (n_10865, n11367);
  and g21592 (n11368, n1296, n_10865);
  not g21593 (n_10866, n11368);
  and g21594 (n11369, n1300, n_10866);
  not g21595 (n_10867, n11369);
  and g21596 (n11370, n1304, n_10867);
  not g21597 (n_10868, n11370);
  and g21598 (n11371, n1308, n_10868);
  not g21599 (n_10869, n11371);
  and g21600 (n11372, n1312, n_10869);
  not g21601 (n_10870, n11372);
  and g21602 (n11373, n1316, n_10870);
  not g21603 (n_10871, n11373);
  and g21604 (n11374, n1320, n_10871);
  not g21605 (n_10872, n11374);
  and g21606 (n11375, n1324, n_10872);
  not g21607 (n_10873, n11375);
  and g21608 (n11376, n1328, n_10873);
  not g21609 (n_10874, n11376);
  and g21610 (n11377, n1332, n_10874);
  not g21611 (n_10875, n11377);
  and g21612 (n11378, n1336, n_10875);
  not g21613 (n_10876, n11378);
  and g21614 (n11379, n1340, n_10876);
  not g21615 (n_10877, n11379);
  and g21616 (n11380, n1344, n_10877);
  not g21617 (n_10878, n11380);
  and g21618 (n11381, n1348, n_10878);
  not g21619 (n_10879, n11381);
  and g21620 (n11382, n1352, n_10879);
  not g21621 (n_10880, n11382);
  and g21622 (n11383, n1356, n_10880);
  not g21623 (n_10881, n11383);
  and g21624 (n11384, n1360, n_10881);
  not g21625 (n_10882, n11384);
  and g21626 (n11385, n1364, n_10882);
  and g21627 (n11386, \req[118] , n_1003);
  not g21628 (n_10883, n11385);
  and g21629 (\grant[118] , n_10883, n11386);
  not g21630 (n_10884, n703);
  and g21631 (n11388, n_10884, n1375);
  not g21632 (n_10885, n11388);
  and g21633 (n11389, n1380, n_10885);
  not g21634 (n_10886, n11389);
  and g21635 (n11390, n1384, n_10886);
  not g21636 (n_10887, n11390);
  and g21637 (n11391, n1388, n_10887);
  not g21638 (n_10888, n11391);
  and g21639 (n11392, n1392, n_10888);
  not g21640 (n_10889, n11392);
  and g21641 (n11393, n1396, n_10889);
  not g21642 (n_10890, n11393);
  and g21643 (n11394, n1663, n_10890);
  not g21644 (n_10891, n11394);
  and g21645 (n11395, n392, n_10891);
  not g21646 (n_10892, n11395);
  and g21647 (n11396, n396, n_10892);
  not g21648 (n_10893, n11396);
  and g21649 (n11397, n400, n_10893);
  not g21650 (n_10894, n11397);
  and g21651 (n11398, n404, n_10894);
  not g21652 (n_10895, n11398);
  and g21653 (n11399, n408, n_10895);
  not g21654 (n_10896, n11399);
  and g21655 (n11400, n412, n_10896);
  not g21656 (n_10897, n11400);
  and g21657 (n11401, n416, n_10897);
  not g21658 (n_10898, n11401);
  and g21659 (n11402, n420, n_10898);
  not g21660 (n_10899, n11402);
  and g21661 (n11403, n424, n_10899);
  not g21662 (n_10900, n11403);
  and g21663 (n11404, n428, n_10900);
  not g21664 (n_10901, n11404);
  and g21665 (n11405, n432, n_10901);
  not g21666 (n_10902, n11405);
  and g21667 (n11406, n436, n_10902);
  not g21668 (n_10903, n11406);
  and g21669 (n11407, n440, n_10903);
  not g21670 (n_10904, n11407);
  and g21671 (n11408, n444, n_10904);
  not g21672 (n_10905, n11408);
  and g21673 (n11409, n448, n_10905);
  not g21674 (n_10906, n11409);
  and g21675 (n11410, n452, n_10906);
  not g21676 (n_10907, n11410);
  and g21677 (n11411, n456, n_10907);
  not g21678 (n_10908, n11411);
  and g21679 (n11412, n460, n_10908);
  not g21680 (n_10909, n11412);
  and g21681 (n11413, n464, n_10909);
  not g21682 (n_10910, n11413);
  and g21683 (n11414, n468, n_10910);
  not g21684 (n_10911, n11414);
  and g21685 (n11415, n472, n_10911);
  not g21686 (n_10912, n11415);
  and g21687 (n11416, n476, n_10912);
  not g21688 (n_10913, n11416);
  and g21689 (n11417, n480, n_10913);
  not g21690 (n_10914, n11417);
  and g21691 (n11418, n484, n_10914);
  not g21692 (n_10915, n11418);
  and g21693 (n11419, n488, n_10915);
  not g21694 (n_10916, n11419);
  and g21695 (n11420, n492, n_10916);
  not g21696 (n_10917, n11420);
  and g21697 (n11421, n496, n_10917);
  not g21698 (n_10918, n11421);
  and g21699 (n11422, n500, n_10918);
  not g21700 (n_10919, n11422);
  and g21701 (n11423, n504, n_10919);
  not g21702 (n_10920, n11423);
  and g21703 (n11424, n508, n_10920);
  not g21704 (n_10921, n11424);
  and g21705 (n11425, n512, n_10921);
  not g21706 (n_10922, n11425);
  and g21707 (n11426, n516, n_10922);
  not g21708 (n_10923, n11426);
  and g21709 (n11427, n520, n_10923);
  not g21710 (n_10924, n11427);
  and g21711 (n11428, n524, n_10924);
  not g21712 (n_10925, n11428);
  and g21713 (n11429, n528, n_10925);
  not g21714 (n_10926, n11429);
  and g21715 (n11430, n532, n_10926);
  not g21716 (n_10927, n11430);
  and g21717 (n11431, n536, n_10927);
  not g21718 (n_10928, n11431);
  and g21719 (n11432, n540, n_10928);
  not g21720 (n_10929, n11432);
  and g21721 (n11433, n544, n_10929);
  not g21722 (n_10930, n11433);
  and g21723 (n11434, n548, n_10930);
  not g21724 (n_10931, n11434);
  and g21725 (n11435, n552, n_10931);
  not g21726 (n_10932, n11435);
  and g21727 (n11436, n556, n_10932);
  not g21728 (n_10933, n11436);
  and g21729 (n11437, n560, n_10933);
  not g21730 (n_10934, n11437);
  and g21731 (n11438, n564, n_10934);
  not g21732 (n_10935, n11438);
  and g21733 (n11439, n568, n_10935);
  not g21734 (n_10936, n11439);
  and g21735 (n11440, n572, n_10936);
  not g21736 (n_10937, n11440);
  and g21737 (n11441, n576, n_10937);
  not g21738 (n_10938, n11441);
  and g21739 (n11442, n580, n_10938);
  not g21740 (n_10939, n11442);
  and g21741 (n11443, n584, n_10939);
  not g21742 (n_10940, n11443);
  and g21743 (n11444, n588, n_10940);
  not g21744 (n_10941, n11444);
  and g21745 (n11445, n592, n_10941);
  not g21746 (n_10942, n11445);
  and g21747 (n11446, n596, n_10942);
  not g21748 (n_10943, n11446);
  and g21749 (n11447, n600, n_10943);
  not g21750 (n_10944, n11447);
  and g21751 (n11448, n604, n_10944);
  not g21752 (n_10945, n11448);
  and g21753 (n11449, n608, n_10945);
  not g21754 (n_10946, n11449);
  and g21755 (n11450, n612, n_10946);
  not g21756 (n_10947, n11450);
  and g21757 (n11451, n616, n_10947);
  not g21758 (n_10948, n11451);
  and g21759 (n11452, n620, n_10948);
  not g21760 (n_10949, n11452);
  and g21761 (n11453, n624, n_10949);
  not g21762 (n_10950, n11453);
  and g21763 (n11454, n628, n_10950);
  not g21764 (n_10951, n11454);
  and g21765 (n11455, n632, n_10951);
  not g21766 (n_10952, n11455);
  and g21767 (n11456, n636, n_10952);
  not g21768 (n_10953, n11456);
  and g21769 (n11457, n640, n_10953);
  not g21770 (n_10954, n11457);
  and g21771 (n11458, n644, n_10954);
  not g21772 (n_10955, n11458);
  and g21773 (n11459, n648, n_10955);
  not g21774 (n_10956, n11459);
  and g21775 (n11460, n652, n_10956);
  not g21776 (n_10957, n11460);
  and g21777 (n11461, n656, n_10957);
  not g21778 (n_10958, n11461);
  and g21779 (n11462, n660, n_10958);
  not g21780 (n_10959, n11462);
  and g21781 (n11463, n664, n_10959);
  not g21782 (n_10960, n11463);
  and g21783 (n11464, n668, n_10960);
  not g21784 (n_10961, n11464);
  and g21785 (n11465, n672, n_10961);
  not g21786 (n_10962, n11465);
  and g21787 (n11466, n676, n_10962);
  not g21788 (n_10963, n11466);
  and g21789 (n11467, n680, n_10963);
  not g21790 (n_10964, n11467);
  and g21791 (n11468, n684, n_10964);
  not g21792 (n_10965, n11468);
  and g21793 (n11469, n688, n_10965);
  not g21794 (n_10966, n11469);
  and g21795 (n11470, n692, n_10966);
  not g21796 (n_10967, n11470);
  and g21797 (n11471, n696, n_10967);
  and g21798 (n11472, \req[119] , n_556);
  not g21799 (n_10968, n11471);
  and g21800 (\grant[119] , n_10968, n11472);
  not g21801 (n_10969, n1042);
  and g21802 (n11474, n707, n_10969);
  not g21803 (n_10970, n11474);
  and g21804 (n11475, n712, n_10970);
  not g21805 (n_10971, n11475);
  and g21806 (n11476, n716, n_10971);
  not g21807 (n_10972, n11476);
  and g21808 (n11477, n720, n_10972);
  not g21809 (n_10973, n11477);
  and g21810 (n11478, n1484, n_10973);
  not g21811 (n_10974, n11478);
  and g21812 (n11479, n1486, n_10974);
  not g21813 (n_10975, n11479);
  and g21814 (n11480, n1750, n_10975);
  not g21815 (n_10976, n11480);
  and g21816 (n11481, n731, n_10976);
  not g21817 (n_10977, n11481);
  and g21818 (n11482, n735, n_10977);
  not g21819 (n_10978, n11482);
  and g21820 (n11483, n739, n_10978);
  not g21821 (n_10979, n11483);
  and g21822 (n11484, n743, n_10979);
  not g21823 (n_10980, n11484);
  and g21824 (n11485, n747, n_10980);
  not g21825 (n_10981, n11485);
  and g21826 (n11486, n751, n_10981);
  not g21827 (n_10982, n11486);
  and g21828 (n11487, n755, n_10982);
  not g21829 (n_10983, n11487);
  and g21830 (n11488, n759, n_10983);
  not g21831 (n_10984, n11488);
  and g21832 (n11489, n763, n_10984);
  not g21833 (n_10985, n11489);
  and g21834 (n11490, n767, n_10985);
  not g21835 (n_10986, n11490);
  and g21836 (n11491, n771, n_10986);
  not g21837 (n_10987, n11491);
  and g21838 (n11492, n775, n_10987);
  not g21839 (n_10988, n11492);
  and g21840 (n11493, n779, n_10988);
  not g21841 (n_10989, n11493);
  and g21842 (n11494, n783, n_10989);
  not g21843 (n_10990, n11494);
  and g21844 (n11495, n787, n_10990);
  not g21845 (n_10991, n11495);
  and g21846 (n11496, n791, n_10991);
  not g21847 (n_10992, n11496);
  and g21848 (n11497, n795, n_10992);
  not g21849 (n_10993, n11497);
  and g21850 (n11498, n799, n_10993);
  not g21851 (n_10994, n11498);
  and g21852 (n11499, n803, n_10994);
  not g21853 (n_10995, n11499);
  and g21854 (n11500, n807, n_10995);
  not g21855 (n_10996, n11500);
  and g21856 (n11501, n811, n_10996);
  not g21857 (n_10997, n11501);
  and g21858 (n11502, n815, n_10997);
  not g21859 (n_10998, n11502);
  and g21860 (n11503, n819, n_10998);
  not g21861 (n_10999, n11503);
  and g21862 (n11504, n823, n_10999);
  not g21863 (n_11000, n11504);
  and g21864 (n11505, n827, n_11000);
  not g21865 (n_11001, n11505);
  and g21866 (n11506, n831, n_11001);
  not g21867 (n_11002, n11506);
  and g21868 (n11507, n835, n_11002);
  not g21869 (n_11003, n11507);
  and g21870 (n11508, n839, n_11003);
  not g21871 (n_11004, n11508);
  and g21872 (n11509, n843, n_11004);
  not g21873 (n_11005, n11509);
  and g21874 (n11510, n847, n_11005);
  not g21875 (n_11006, n11510);
  and g21876 (n11511, n851, n_11006);
  not g21877 (n_11007, n11511);
  and g21878 (n11512, n855, n_11007);
  not g21879 (n_11008, n11512);
  and g21880 (n11513, n859, n_11008);
  not g21881 (n_11009, n11513);
  and g21882 (n11514, n863, n_11009);
  not g21883 (n_11010, n11514);
  and g21884 (n11515, n867, n_11010);
  not g21885 (n_11011, n11515);
  and g21886 (n11516, n871, n_11011);
  not g21887 (n_11012, n11516);
  and g21888 (n11517, n875, n_11012);
  not g21889 (n_11013, n11517);
  and g21890 (n11518, n879, n_11013);
  not g21891 (n_11014, n11518);
  and g21892 (n11519, n883, n_11014);
  not g21893 (n_11015, n11519);
  and g21894 (n11520, n887, n_11015);
  not g21895 (n_11016, n11520);
  and g21896 (n11521, n891, n_11016);
  not g21897 (n_11017, n11521);
  and g21898 (n11522, n895, n_11017);
  not g21899 (n_11018, n11522);
  and g21900 (n11523, n899, n_11018);
  not g21901 (n_11019, n11523);
  and g21902 (n11524, n903, n_11019);
  not g21903 (n_11020, n11524);
  and g21904 (n11525, n907, n_11020);
  not g21905 (n_11021, n11525);
  and g21906 (n11526, n911, n_11021);
  not g21907 (n_11022, n11526);
  and g21908 (n11527, n915, n_11022);
  not g21909 (n_11023, n11527);
  and g21910 (n11528, n919, n_11023);
  not g21911 (n_11024, n11528);
  and g21912 (n11529, n923, n_11024);
  not g21913 (n_11025, n11529);
  and g21914 (n11530, n927, n_11025);
  not g21915 (n_11026, n11530);
  and g21916 (n11531, n931, n_11026);
  not g21917 (n_11027, n11531);
  and g21918 (n11532, n935, n_11027);
  not g21919 (n_11028, n11532);
  and g21920 (n11533, n939, n_11028);
  not g21921 (n_11029, n11533);
  and g21922 (n11534, n943, n_11029);
  not g21923 (n_11030, n11534);
  and g21924 (n11535, n947, n_11030);
  not g21925 (n_11031, n11535);
  and g21926 (n11536, n951, n_11031);
  not g21927 (n_11032, n11536);
  and g21928 (n11537, n955, n_11032);
  not g21929 (n_11033, n11537);
  and g21930 (n11538, n959, n_11033);
  not g21931 (n_11034, n11538);
  and g21932 (n11539, n963, n_11034);
  not g21933 (n_11035, n11539);
  and g21934 (n11540, n967, n_11035);
  not g21935 (n_11036, n11540);
  and g21936 (n11541, n971, n_11036);
  not g21937 (n_11037, n11541);
  and g21938 (n11542, n975, n_11037);
  not g21939 (n_11038, n11542);
  and g21940 (n11543, n979, n_11038);
  not g21941 (n_11039, n11543);
  and g21942 (n11544, n983, n_11039);
  not g21943 (n_11040, n11544);
  and g21944 (n11545, n987, n_11040);
  not g21945 (n_11041, n11545);
  and g21946 (n11546, n991, n_11041);
  not g21947 (n_11042, n11546);
  and g21948 (n11547, n995, n_11042);
  not g21949 (n_11043, n11547);
  and g21950 (n11548, n999, n_11043);
  not g21951 (n_11044, n11548);
  and g21952 (n11549, n1003, n_11044);
  not g21953 (n_11045, n11549);
  and g21954 (n11550, n1007, n_11045);
  not g21955 (n_11046, n11550);
  and g21956 (n11551, n1011, n_11046);
  not g21957 (n_11047, n11551);
  and g21958 (n11552, n1015, n_11047);
  not g21959 (n_11048, n11552);
  and g21960 (n11553, n1019, n_11048);
  not g21961 (n_11049, n11553);
  and g21962 (n11554, n1023, n_11049);
  not g21963 (n_11050, n11554);
  and g21964 (n11555, n1027, n_11050);
  not g21965 (n_11051, n11555);
  and g21966 (n11556, n1031, n_11051);
  not g21967 (n_11052, n11556);
  and g21968 (n11557, n1035, n_11052);
  and g21969 (n11558, \req[120] , n_833);
  not g21970 (n_11053, n11557);
  and g21971 (\grant[120] , n_11053, n11558);
  not g21972 (n_11054, n1379);
  and g21973 (n11560, n1046, n_11054);
  not g21974 (n_11055, n11560);
  and g21975 (n11561, n1051, n_11055);
  not g21976 (n_11056, n11561);
  and g21977 (n11562, n1055, n_11056);
  not g21978 (n_11057, n11562);
  and g21979 (n11563, n1059, n_11057);
  not g21980 (n_11058, n11563);
  and g21981 (n11564, n1574, n_11058);
  not g21982 (n_11059, n11564);
  and g21983 (n11565, n1576, n_11059);
  not g21984 (n_11060, n11565);
  and g21985 (n11566, n1837, n_11060);
  not g21986 (n_11061, n11566);
  and g21987 (n11567, n1068, n_11061);
  not g21988 (n_11062, n11567);
  and g21989 (n11568, n1072, n_11062);
  not g21990 (n_11063, n11568);
  and g21991 (n11569, n1076, n_11063);
  not g21992 (n_11064, n11569);
  and g21993 (n11570, n1080, n_11064);
  not g21994 (n_11065, n11570);
  and g21995 (n11571, n1084, n_11065);
  not g21996 (n_11066, n11571);
  and g21997 (n11572, n1088, n_11066);
  not g21998 (n_11067, n11572);
  and g21999 (n11573, n1092, n_11067);
  not g22000 (n_11068, n11573);
  and g22001 (n11574, n1096, n_11068);
  not g22002 (n_11069, n11574);
  and g22003 (n11575, n1100, n_11069);
  not g22004 (n_11070, n11575);
  and g22005 (n11576, n1104, n_11070);
  not g22006 (n_11071, n11576);
  and g22007 (n11577, n1108, n_11071);
  not g22008 (n_11072, n11577);
  and g22009 (n11578, n1112, n_11072);
  not g22010 (n_11073, n11578);
  and g22011 (n11579, n1116, n_11073);
  not g22012 (n_11074, n11579);
  and g22013 (n11580, n1120, n_11074);
  not g22014 (n_11075, n11580);
  and g22015 (n11581, n1124, n_11075);
  not g22016 (n_11076, n11581);
  and g22017 (n11582, n1128, n_11076);
  not g22018 (n_11077, n11582);
  and g22019 (n11583, n1132, n_11077);
  not g22020 (n_11078, n11583);
  and g22021 (n11584, n1136, n_11078);
  not g22022 (n_11079, n11584);
  and g22023 (n11585, n1140, n_11079);
  not g22024 (n_11080, n11585);
  and g22025 (n11586, n1144, n_11080);
  not g22026 (n_11081, n11586);
  and g22027 (n11587, n1148, n_11081);
  not g22028 (n_11082, n11587);
  and g22029 (n11588, n1152, n_11082);
  not g22030 (n_11083, n11588);
  and g22031 (n11589, n1156, n_11083);
  not g22032 (n_11084, n11589);
  and g22033 (n11590, n1160, n_11084);
  not g22034 (n_11085, n11590);
  and g22035 (n11591, n1164, n_11085);
  not g22036 (n_11086, n11591);
  and g22037 (n11592, n1168, n_11086);
  not g22038 (n_11087, n11592);
  and g22039 (n11593, n1172, n_11087);
  not g22040 (n_11088, n11593);
  and g22041 (n11594, n1176, n_11088);
  not g22042 (n_11089, n11594);
  and g22043 (n11595, n1180, n_11089);
  not g22044 (n_11090, n11595);
  and g22045 (n11596, n1184, n_11090);
  not g22046 (n_11091, n11596);
  and g22047 (n11597, n1188, n_11091);
  not g22048 (n_11092, n11597);
  and g22049 (n11598, n1192, n_11092);
  not g22050 (n_11093, n11598);
  and g22051 (n11599, n1196, n_11093);
  not g22052 (n_11094, n11599);
  and g22053 (n11600, n1200, n_11094);
  not g22054 (n_11095, n11600);
  and g22055 (n11601, n1204, n_11095);
  not g22056 (n_11096, n11601);
  and g22057 (n11602, n1208, n_11096);
  not g22058 (n_11097, n11602);
  and g22059 (n11603, n1212, n_11097);
  not g22060 (n_11098, n11603);
  and g22061 (n11604, n1216, n_11098);
  not g22062 (n_11099, n11604);
  and g22063 (n11605, n1220, n_11099);
  not g22064 (n_11100, n11605);
  and g22065 (n11606, n1224, n_11100);
  not g22066 (n_11101, n11606);
  and g22067 (n11607, n1228, n_11101);
  not g22068 (n_11102, n11607);
  and g22069 (n11608, n1232, n_11102);
  not g22070 (n_11103, n11608);
  and g22071 (n11609, n1236, n_11103);
  not g22072 (n_11104, n11609);
  and g22073 (n11610, n1240, n_11104);
  not g22074 (n_11105, n11610);
  and g22075 (n11611, n1244, n_11105);
  not g22076 (n_11106, n11611);
  and g22077 (n11612, n1248, n_11106);
  not g22078 (n_11107, n11612);
  and g22079 (n11613, n1252, n_11107);
  not g22080 (n_11108, n11613);
  and g22081 (n11614, n1256, n_11108);
  not g22082 (n_11109, n11614);
  and g22083 (n11615, n1260, n_11109);
  not g22084 (n_11110, n11615);
  and g22085 (n11616, n1264, n_11110);
  not g22086 (n_11111, n11616);
  and g22087 (n11617, n1268, n_11111);
  not g22088 (n_11112, n11617);
  and g22089 (n11618, n1272, n_11112);
  not g22090 (n_11113, n11618);
  and g22091 (n11619, n1276, n_11113);
  not g22092 (n_11114, n11619);
  and g22093 (n11620, n1280, n_11114);
  not g22094 (n_11115, n11620);
  and g22095 (n11621, n1284, n_11115);
  not g22096 (n_11116, n11621);
  and g22097 (n11622, n1288, n_11116);
  not g22098 (n_11117, n11622);
  and g22099 (n11623, n1292, n_11117);
  not g22100 (n_11118, n11623);
  and g22101 (n11624, n1296, n_11118);
  not g22102 (n_11119, n11624);
  and g22103 (n11625, n1300, n_11119);
  not g22104 (n_11120, n11625);
  and g22105 (n11626, n1304, n_11120);
  not g22106 (n_11121, n11626);
  and g22107 (n11627, n1308, n_11121);
  not g22108 (n_11122, n11627);
  and g22109 (n11628, n1312, n_11122);
  not g22110 (n_11123, n11628);
  and g22111 (n11629, n1316, n_11123);
  not g22112 (n_11124, n11629);
  and g22113 (n11630, n1320, n_11124);
  not g22114 (n_11125, n11630);
  and g22115 (n11631, n1324, n_11125);
  not g22116 (n_11126, n11631);
  and g22117 (n11632, n1328, n_11126);
  not g22118 (n_11127, n11632);
  and g22119 (n11633, n1332, n_11127);
  not g22120 (n_11128, n11633);
  and g22121 (n11634, n1336, n_11128);
  not g22122 (n_11129, n11634);
  and g22123 (n11635, n1340, n_11129);
  not g22124 (n_11130, n11635);
  and g22125 (n11636, n1344, n_11130);
  not g22126 (n_11131, n11636);
  and g22127 (n11637, n1348, n_11131);
  not g22128 (n_11132, n11637);
  and g22129 (n11638, n1352, n_11132);
  not g22130 (n_11133, n11638);
  and g22131 (n11639, n1356, n_11133);
  not g22132 (n_11134, n11639);
  and g22133 (n11640, n1360, n_11134);
  not g22134 (n_11135, n11640);
  and g22135 (n11641, n1364, n_11135);
  not g22136 (n_11136, n11641);
  and g22137 (n11642, n1368, n_11136);
  not g22138 (n_11137, n11642);
  and g22139 (n11643, n1372, n_11137);
  and g22140 (n11644, \req[121] , n_1007);
  not g22141 (n_11138, n11643);
  and g22142 (\grant[121] , n_11138, n11644);
  not g22143 (n_11139, n711);
  and g22144 (n11646, n_11139, n1383);
  not g22145 (n_11140, n11646);
  and g22146 (n11647, n1388, n_11140);
  not g22147 (n_11141, n11647);
  and g22148 (n11648, n1392, n_11141);
  not g22149 (n_11142, n11648);
  and g22150 (n11649, n1396, n_11142);
  not g22151 (n_11143, n11649);
  and g22152 (n11650, n1663, n_11143);
  not g22153 (n_11144, n11650);
  and g22154 (n11651, n392, n_11144);
  not g22155 (n_11145, n11651);
  and g22156 (n11652, n396, n_11145);
  not g22157 (n_11146, n11652);
  and g22158 (n11653, n400, n_11146);
  not g22159 (n_11147, n11653);
  and g22160 (n11654, n404, n_11147);
  not g22161 (n_11148, n11654);
  and g22162 (n11655, n408, n_11148);
  not g22163 (n_11149, n11655);
  and g22164 (n11656, n412, n_11149);
  not g22165 (n_11150, n11656);
  and g22166 (n11657, n416, n_11150);
  not g22167 (n_11151, n11657);
  and g22168 (n11658, n420, n_11151);
  not g22169 (n_11152, n11658);
  and g22170 (n11659, n424, n_11152);
  not g22171 (n_11153, n11659);
  and g22172 (n11660, n428, n_11153);
  not g22173 (n_11154, n11660);
  and g22174 (n11661, n432, n_11154);
  not g22175 (n_11155, n11661);
  and g22176 (n11662, n436, n_11155);
  not g22177 (n_11156, n11662);
  and g22178 (n11663, n440, n_11156);
  not g22179 (n_11157, n11663);
  and g22180 (n11664, n444, n_11157);
  not g22181 (n_11158, n11664);
  and g22182 (n11665, n448, n_11158);
  not g22183 (n_11159, n11665);
  and g22184 (n11666, n452, n_11159);
  not g22185 (n_11160, n11666);
  and g22186 (n11667, n456, n_11160);
  not g22187 (n_11161, n11667);
  and g22188 (n11668, n460, n_11161);
  not g22189 (n_11162, n11668);
  and g22190 (n11669, n464, n_11162);
  not g22191 (n_11163, n11669);
  and g22192 (n11670, n468, n_11163);
  not g22193 (n_11164, n11670);
  and g22194 (n11671, n472, n_11164);
  not g22195 (n_11165, n11671);
  and g22196 (n11672, n476, n_11165);
  not g22197 (n_11166, n11672);
  and g22198 (n11673, n480, n_11166);
  not g22199 (n_11167, n11673);
  and g22200 (n11674, n484, n_11167);
  not g22201 (n_11168, n11674);
  and g22202 (n11675, n488, n_11168);
  not g22203 (n_11169, n11675);
  and g22204 (n11676, n492, n_11169);
  not g22205 (n_11170, n11676);
  and g22206 (n11677, n496, n_11170);
  not g22207 (n_11171, n11677);
  and g22208 (n11678, n500, n_11171);
  not g22209 (n_11172, n11678);
  and g22210 (n11679, n504, n_11172);
  not g22211 (n_11173, n11679);
  and g22212 (n11680, n508, n_11173);
  not g22213 (n_11174, n11680);
  and g22214 (n11681, n512, n_11174);
  not g22215 (n_11175, n11681);
  and g22216 (n11682, n516, n_11175);
  not g22217 (n_11176, n11682);
  and g22218 (n11683, n520, n_11176);
  not g22219 (n_11177, n11683);
  and g22220 (n11684, n524, n_11177);
  not g22221 (n_11178, n11684);
  and g22222 (n11685, n528, n_11178);
  not g22223 (n_11179, n11685);
  and g22224 (n11686, n532, n_11179);
  not g22225 (n_11180, n11686);
  and g22226 (n11687, n536, n_11180);
  not g22227 (n_11181, n11687);
  and g22228 (n11688, n540, n_11181);
  not g22229 (n_11182, n11688);
  and g22230 (n11689, n544, n_11182);
  not g22231 (n_11183, n11689);
  and g22232 (n11690, n548, n_11183);
  not g22233 (n_11184, n11690);
  and g22234 (n11691, n552, n_11184);
  not g22235 (n_11185, n11691);
  and g22236 (n11692, n556, n_11185);
  not g22237 (n_11186, n11692);
  and g22238 (n11693, n560, n_11186);
  not g22239 (n_11187, n11693);
  and g22240 (n11694, n564, n_11187);
  not g22241 (n_11188, n11694);
  and g22242 (n11695, n568, n_11188);
  not g22243 (n_11189, n11695);
  and g22244 (n11696, n572, n_11189);
  not g22245 (n_11190, n11696);
  and g22246 (n11697, n576, n_11190);
  not g22247 (n_11191, n11697);
  and g22248 (n11698, n580, n_11191);
  not g22249 (n_11192, n11698);
  and g22250 (n11699, n584, n_11192);
  not g22251 (n_11193, n11699);
  and g22252 (n11700, n588, n_11193);
  not g22253 (n_11194, n11700);
  and g22254 (n11701, n592, n_11194);
  not g22255 (n_11195, n11701);
  and g22256 (n11702, n596, n_11195);
  not g22257 (n_11196, n11702);
  and g22258 (n11703, n600, n_11196);
  not g22259 (n_11197, n11703);
  and g22260 (n11704, n604, n_11197);
  not g22261 (n_11198, n11704);
  and g22262 (n11705, n608, n_11198);
  not g22263 (n_11199, n11705);
  and g22264 (n11706, n612, n_11199);
  not g22265 (n_11200, n11706);
  and g22266 (n11707, n616, n_11200);
  not g22267 (n_11201, n11707);
  and g22268 (n11708, n620, n_11201);
  not g22269 (n_11202, n11708);
  and g22270 (n11709, n624, n_11202);
  not g22271 (n_11203, n11709);
  and g22272 (n11710, n628, n_11203);
  not g22273 (n_11204, n11710);
  and g22274 (n11711, n632, n_11204);
  not g22275 (n_11205, n11711);
  and g22276 (n11712, n636, n_11205);
  not g22277 (n_11206, n11712);
  and g22278 (n11713, n640, n_11206);
  not g22279 (n_11207, n11713);
  and g22280 (n11714, n644, n_11207);
  not g22281 (n_11208, n11714);
  and g22282 (n11715, n648, n_11208);
  not g22283 (n_11209, n11715);
  and g22284 (n11716, n652, n_11209);
  not g22285 (n_11210, n11716);
  and g22286 (n11717, n656, n_11210);
  not g22287 (n_11211, n11717);
  and g22288 (n11718, n660, n_11211);
  not g22289 (n_11212, n11718);
  and g22290 (n11719, n664, n_11212);
  not g22291 (n_11213, n11719);
  and g22292 (n11720, n668, n_11213);
  not g22293 (n_11214, n11720);
  and g22294 (n11721, n672, n_11214);
  not g22295 (n_11215, n11721);
  and g22296 (n11722, n676, n_11215);
  not g22297 (n_11216, n11722);
  and g22298 (n11723, n680, n_11216);
  not g22299 (n_11217, n11723);
  and g22300 (n11724, n684, n_11217);
  not g22301 (n_11218, n11724);
  and g22302 (n11725, n688, n_11218);
  not g22303 (n_11219, n11725);
  and g22304 (n11726, n692, n_11219);
  not g22305 (n_11220, n11726);
  and g22306 (n11727, n696, n_11220);
  not g22307 (n_11221, n11727);
  and g22308 (n11728, n700, n_11221);
  not g22309 (n_11222, n11728);
  and g22310 (n11729, n704, n_11222);
  and g22311 (n11730, \req[122] , n_570);
  not g22312 (n_11223, n11729);
  and g22313 (\grant[122] , n_11223, n11730);
  not g22314 (n_11224, n1050);
  and g22315 (n11732, n715, n_11224);
  not g22316 (n_11225, n11732);
  and g22317 (n11733, n720, n_11225);
  not g22318 (n_11226, n11733);
  and g22319 (n11734, n1484, n_11226);
  not g22320 (n_11227, n11734);
  and g22321 (n11735, n1486, n_11227);
  not g22322 (n_11228, n11735);
  and g22323 (n11736, n1750, n_11228);
  not g22324 (n_11229, n11736);
  and g22325 (n11737, n731, n_11229);
  not g22326 (n_11230, n11737);
  and g22327 (n11738, n735, n_11230);
  not g22328 (n_11231, n11738);
  and g22329 (n11739, n739, n_11231);
  not g22330 (n_11232, n11739);
  and g22331 (n11740, n743, n_11232);
  not g22332 (n_11233, n11740);
  and g22333 (n11741, n747, n_11233);
  not g22334 (n_11234, n11741);
  and g22335 (n11742, n751, n_11234);
  not g22336 (n_11235, n11742);
  and g22337 (n11743, n755, n_11235);
  not g22338 (n_11236, n11743);
  and g22339 (n11744, n759, n_11236);
  not g22340 (n_11237, n11744);
  and g22341 (n11745, n763, n_11237);
  not g22342 (n_11238, n11745);
  and g22343 (n11746, n767, n_11238);
  not g22344 (n_11239, n11746);
  and g22345 (n11747, n771, n_11239);
  not g22346 (n_11240, n11747);
  and g22347 (n11748, n775, n_11240);
  not g22348 (n_11241, n11748);
  and g22349 (n11749, n779, n_11241);
  not g22350 (n_11242, n11749);
  and g22351 (n11750, n783, n_11242);
  not g22352 (n_11243, n11750);
  and g22353 (n11751, n787, n_11243);
  not g22354 (n_11244, n11751);
  and g22355 (n11752, n791, n_11244);
  not g22356 (n_11245, n11752);
  and g22357 (n11753, n795, n_11245);
  not g22358 (n_11246, n11753);
  and g22359 (n11754, n799, n_11246);
  not g22360 (n_11247, n11754);
  and g22361 (n11755, n803, n_11247);
  not g22362 (n_11248, n11755);
  and g22363 (n11756, n807, n_11248);
  not g22364 (n_11249, n11756);
  and g22365 (n11757, n811, n_11249);
  not g22366 (n_11250, n11757);
  and g22367 (n11758, n815, n_11250);
  not g22368 (n_11251, n11758);
  and g22369 (n11759, n819, n_11251);
  not g22370 (n_11252, n11759);
  and g22371 (n11760, n823, n_11252);
  not g22372 (n_11253, n11760);
  and g22373 (n11761, n827, n_11253);
  not g22374 (n_11254, n11761);
  and g22375 (n11762, n831, n_11254);
  not g22376 (n_11255, n11762);
  and g22377 (n11763, n835, n_11255);
  not g22378 (n_11256, n11763);
  and g22379 (n11764, n839, n_11256);
  not g22380 (n_11257, n11764);
  and g22381 (n11765, n843, n_11257);
  not g22382 (n_11258, n11765);
  and g22383 (n11766, n847, n_11258);
  not g22384 (n_11259, n11766);
  and g22385 (n11767, n851, n_11259);
  not g22386 (n_11260, n11767);
  and g22387 (n11768, n855, n_11260);
  not g22388 (n_11261, n11768);
  and g22389 (n11769, n859, n_11261);
  not g22390 (n_11262, n11769);
  and g22391 (n11770, n863, n_11262);
  not g22392 (n_11263, n11770);
  and g22393 (n11771, n867, n_11263);
  not g22394 (n_11264, n11771);
  and g22395 (n11772, n871, n_11264);
  not g22396 (n_11265, n11772);
  and g22397 (n11773, n875, n_11265);
  not g22398 (n_11266, n11773);
  and g22399 (n11774, n879, n_11266);
  not g22400 (n_11267, n11774);
  and g22401 (n11775, n883, n_11267);
  not g22402 (n_11268, n11775);
  and g22403 (n11776, n887, n_11268);
  not g22404 (n_11269, n11776);
  and g22405 (n11777, n891, n_11269);
  not g22406 (n_11270, n11777);
  and g22407 (n11778, n895, n_11270);
  not g22408 (n_11271, n11778);
  and g22409 (n11779, n899, n_11271);
  not g22410 (n_11272, n11779);
  and g22411 (n11780, n903, n_11272);
  not g22412 (n_11273, n11780);
  and g22413 (n11781, n907, n_11273);
  not g22414 (n_11274, n11781);
  and g22415 (n11782, n911, n_11274);
  not g22416 (n_11275, n11782);
  and g22417 (n11783, n915, n_11275);
  not g22418 (n_11276, n11783);
  and g22419 (n11784, n919, n_11276);
  not g22420 (n_11277, n11784);
  and g22421 (n11785, n923, n_11277);
  not g22422 (n_11278, n11785);
  and g22423 (n11786, n927, n_11278);
  not g22424 (n_11279, n11786);
  and g22425 (n11787, n931, n_11279);
  not g22426 (n_11280, n11787);
  and g22427 (n11788, n935, n_11280);
  not g22428 (n_11281, n11788);
  and g22429 (n11789, n939, n_11281);
  not g22430 (n_11282, n11789);
  and g22431 (n11790, n943, n_11282);
  not g22432 (n_11283, n11790);
  and g22433 (n11791, n947, n_11283);
  not g22434 (n_11284, n11791);
  and g22435 (n11792, n951, n_11284);
  not g22436 (n_11285, n11792);
  and g22437 (n11793, n955, n_11285);
  not g22438 (n_11286, n11793);
  and g22439 (n11794, n959, n_11286);
  not g22440 (n_11287, n11794);
  and g22441 (n11795, n963, n_11287);
  not g22442 (n_11288, n11795);
  and g22443 (n11796, n967, n_11288);
  not g22444 (n_11289, n11796);
  and g22445 (n11797, n971, n_11289);
  not g22446 (n_11290, n11797);
  and g22447 (n11798, n975, n_11290);
  not g22448 (n_11291, n11798);
  and g22449 (n11799, n979, n_11291);
  not g22450 (n_11292, n11799);
  and g22451 (n11800, n983, n_11292);
  not g22452 (n_11293, n11800);
  and g22453 (n11801, n987, n_11293);
  not g22454 (n_11294, n11801);
  and g22455 (n11802, n991, n_11294);
  not g22456 (n_11295, n11802);
  and g22457 (n11803, n995, n_11295);
  not g22458 (n_11296, n11803);
  and g22459 (n11804, n999, n_11296);
  not g22460 (n_11297, n11804);
  and g22461 (n11805, n1003, n_11297);
  not g22462 (n_11298, n11805);
  and g22463 (n11806, n1007, n_11298);
  not g22464 (n_11299, n11806);
  and g22465 (n11807, n1011, n_11299);
  not g22466 (n_11300, n11807);
  and g22467 (n11808, n1015, n_11300);
  not g22468 (n_11301, n11808);
  and g22469 (n11809, n1019, n_11301);
  not g22470 (n_11302, n11809);
  and g22471 (n11810, n1023, n_11302);
  not g22472 (n_11303, n11810);
  and g22473 (n11811, n1027, n_11303);
  not g22474 (n_11304, n11811);
  and g22475 (n11812, n1031, n_11304);
  not g22476 (n_11305, n11812);
  and g22477 (n11813, n1035, n_11305);
  not g22478 (n_11306, n11813);
  and g22479 (n11814, n1039, n_11306);
  not g22480 (n_11307, n11814);
  and g22481 (n11815, n1043, n_11307);
  and g22482 (n11816, \req[123] , n_839);
  not g22483 (n_11308, n11815);
  and g22484 (\grant[123] , n_11308, n11816);
  not g22485 (n_11309, n1387);
  and g22486 (n11818, n1054, n_11309);
  not g22487 (n_11310, n11818);
  and g22488 (n11819, n1059, n_11310);
  not g22489 (n_11311, n11819);
  and g22490 (n11820, n1574, n_11311);
  not g22491 (n_11312, n11820);
  and g22492 (n11821, n1576, n_11312);
  not g22493 (n_11313, n11821);
  and g22494 (n11822, n1837, n_11313);
  not g22495 (n_11314, n11822);
  and g22496 (n11823, n1068, n_11314);
  not g22497 (n_11315, n11823);
  and g22498 (n11824, n1072, n_11315);
  not g22499 (n_11316, n11824);
  and g22500 (n11825, n1076, n_11316);
  not g22501 (n_11317, n11825);
  and g22502 (n11826, n1080, n_11317);
  not g22503 (n_11318, n11826);
  and g22504 (n11827, n1084, n_11318);
  not g22505 (n_11319, n11827);
  and g22506 (n11828, n1088, n_11319);
  not g22507 (n_11320, n11828);
  and g22508 (n11829, n1092, n_11320);
  not g22509 (n_11321, n11829);
  and g22510 (n11830, n1096, n_11321);
  not g22511 (n_11322, n11830);
  and g22512 (n11831, n1100, n_11322);
  not g22513 (n_11323, n11831);
  and g22514 (n11832, n1104, n_11323);
  not g22515 (n_11324, n11832);
  and g22516 (n11833, n1108, n_11324);
  not g22517 (n_11325, n11833);
  and g22518 (n11834, n1112, n_11325);
  not g22519 (n_11326, n11834);
  and g22520 (n11835, n1116, n_11326);
  not g22521 (n_11327, n11835);
  and g22522 (n11836, n1120, n_11327);
  not g22523 (n_11328, n11836);
  and g22524 (n11837, n1124, n_11328);
  not g22525 (n_11329, n11837);
  and g22526 (n11838, n1128, n_11329);
  not g22527 (n_11330, n11838);
  and g22528 (n11839, n1132, n_11330);
  not g22529 (n_11331, n11839);
  and g22530 (n11840, n1136, n_11331);
  not g22531 (n_11332, n11840);
  and g22532 (n11841, n1140, n_11332);
  not g22533 (n_11333, n11841);
  and g22534 (n11842, n1144, n_11333);
  not g22535 (n_11334, n11842);
  and g22536 (n11843, n1148, n_11334);
  not g22537 (n_11335, n11843);
  and g22538 (n11844, n1152, n_11335);
  not g22539 (n_11336, n11844);
  and g22540 (n11845, n1156, n_11336);
  not g22541 (n_11337, n11845);
  and g22542 (n11846, n1160, n_11337);
  not g22543 (n_11338, n11846);
  and g22544 (n11847, n1164, n_11338);
  not g22545 (n_11339, n11847);
  and g22546 (n11848, n1168, n_11339);
  not g22547 (n_11340, n11848);
  and g22548 (n11849, n1172, n_11340);
  not g22549 (n_11341, n11849);
  and g22550 (n11850, n1176, n_11341);
  not g22551 (n_11342, n11850);
  and g22552 (n11851, n1180, n_11342);
  not g22553 (n_11343, n11851);
  and g22554 (n11852, n1184, n_11343);
  not g22555 (n_11344, n11852);
  and g22556 (n11853, n1188, n_11344);
  not g22557 (n_11345, n11853);
  and g22558 (n11854, n1192, n_11345);
  not g22559 (n_11346, n11854);
  and g22560 (n11855, n1196, n_11346);
  not g22561 (n_11347, n11855);
  and g22562 (n11856, n1200, n_11347);
  not g22563 (n_11348, n11856);
  and g22564 (n11857, n1204, n_11348);
  not g22565 (n_11349, n11857);
  and g22566 (n11858, n1208, n_11349);
  not g22567 (n_11350, n11858);
  and g22568 (n11859, n1212, n_11350);
  not g22569 (n_11351, n11859);
  and g22570 (n11860, n1216, n_11351);
  not g22571 (n_11352, n11860);
  and g22572 (n11861, n1220, n_11352);
  not g22573 (n_11353, n11861);
  and g22574 (n11862, n1224, n_11353);
  not g22575 (n_11354, n11862);
  and g22576 (n11863, n1228, n_11354);
  not g22577 (n_11355, n11863);
  and g22578 (n11864, n1232, n_11355);
  not g22579 (n_11356, n11864);
  and g22580 (n11865, n1236, n_11356);
  not g22581 (n_11357, n11865);
  and g22582 (n11866, n1240, n_11357);
  not g22583 (n_11358, n11866);
  and g22584 (n11867, n1244, n_11358);
  not g22585 (n_11359, n11867);
  and g22586 (n11868, n1248, n_11359);
  not g22587 (n_11360, n11868);
  and g22588 (n11869, n1252, n_11360);
  not g22589 (n_11361, n11869);
  and g22590 (n11870, n1256, n_11361);
  not g22591 (n_11362, n11870);
  and g22592 (n11871, n1260, n_11362);
  not g22593 (n_11363, n11871);
  and g22594 (n11872, n1264, n_11363);
  not g22595 (n_11364, n11872);
  and g22596 (n11873, n1268, n_11364);
  not g22597 (n_11365, n11873);
  and g22598 (n11874, n1272, n_11365);
  not g22599 (n_11366, n11874);
  and g22600 (n11875, n1276, n_11366);
  not g22601 (n_11367, n11875);
  and g22602 (n11876, n1280, n_11367);
  not g22603 (n_11368, n11876);
  and g22604 (n11877, n1284, n_11368);
  not g22605 (n_11369, n11877);
  and g22606 (n11878, n1288, n_11369);
  not g22607 (n_11370, n11878);
  and g22608 (n11879, n1292, n_11370);
  not g22609 (n_11371, n11879);
  and g22610 (n11880, n1296, n_11371);
  not g22611 (n_11372, n11880);
  and g22612 (n11881, n1300, n_11372);
  not g22613 (n_11373, n11881);
  and g22614 (n11882, n1304, n_11373);
  not g22615 (n_11374, n11882);
  and g22616 (n11883, n1308, n_11374);
  not g22617 (n_11375, n11883);
  and g22618 (n11884, n1312, n_11375);
  not g22619 (n_11376, n11884);
  and g22620 (n11885, n1316, n_11376);
  not g22621 (n_11377, n11885);
  and g22622 (n11886, n1320, n_11377);
  not g22623 (n_11378, n11886);
  and g22624 (n11887, n1324, n_11378);
  not g22625 (n_11379, n11887);
  and g22626 (n11888, n1328, n_11379);
  not g22627 (n_11380, n11888);
  and g22628 (n11889, n1332, n_11380);
  not g22629 (n_11381, n11889);
  and g22630 (n11890, n1336, n_11381);
  not g22631 (n_11382, n11890);
  and g22632 (n11891, n1340, n_11382);
  not g22633 (n_11383, n11891);
  and g22634 (n11892, n1344, n_11383);
  not g22635 (n_11384, n11892);
  and g22636 (n11893, n1348, n_11384);
  not g22637 (n_11385, n11893);
  and g22638 (n11894, n1352, n_11385);
  not g22639 (n_11386, n11894);
  and g22640 (n11895, n1356, n_11386);
  not g22641 (n_11387, n11895);
  and g22642 (n11896, n1360, n_11387);
  not g22643 (n_11388, n11896);
  and g22644 (n11897, n1364, n_11388);
  not g22645 (n_11389, n11897);
  and g22646 (n11898, n1368, n_11389);
  not g22647 (n_11390, n11898);
  and g22648 (n11899, n1372, n_11390);
  not g22649 (n_11391, n11899);
  and g22650 (n11900, n1376, n_11391);
  not g22651 (n_11392, n11900);
  and g22652 (n11901, n1380, n_11392);
  and g22653 (n11902, \req[124] , n_1011);
  not g22654 (n_11393, n11901);
  and g22655 (\grant[124] , n_11393, n11902);
  not g22656 (n_11394, n719);
  and g22657 (n11904, n_11394, n1391);
  not g22658 (n_11395, n11904);
  and g22659 (n11905, n1396, n_11395);
  not g22660 (n_11396, n11905);
  and g22661 (n11906, n1663, n_11396);
  not g22662 (n_11397, n11906);
  and g22663 (n11907, n392, n_11397);
  not g22664 (n_11398, n11907);
  and g22665 (n11908, n396, n_11398);
  not g22666 (n_11399, n11908);
  and g22667 (n11909, n400, n_11399);
  not g22668 (n_11400, n11909);
  and g22669 (n11910, n404, n_11400);
  not g22670 (n_11401, n11910);
  and g22671 (n11911, n408, n_11401);
  not g22672 (n_11402, n11911);
  and g22673 (n11912, n412, n_11402);
  not g22674 (n_11403, n11912);
  and g22675 (n11913, n416, n_11403);
  not g22676 (n_11404, n11913);
  and g22677 (n11914, n420, n_11404);
  not g22678 (n_11405, n11914);
  and g22679 (n11915, n424, n_11405);
  not g22680 (n_11406, n11915);
  and g22681 (n11916, n428, n_11406);
  not g22682 (n_11407, n11916);
  and g22683 (n11917, n432, n_11407);
  not g22684 (n_11408, n11917);
  and g22685 (n11918, n436, n_11408);
  not g22686 (n_11409, n11918);
  and g22687 (n11919, n440, n_11409);
  not g22688 (n_11410, n11919);
  and g22689 (n11920, n444, n_11410);
  not g22690 (n_11411, n11920);
  and g22691 (n11921, n448, n_11411);
  not g22692 (n_11412, n11921);
  and g22693 (n11922, n452, n_11412);
  not g22694 (n_11413, n11922);
  and g22695 (n11923, n456, n_11413);
  not g22696 (n_11414, n11923);
  and g22697 (n11924, n460, n_11414);
  not g22698 (n_11415, n11924);
  and g22699 (n11925, n464, n_11415);
  not g22700 (n_11416, n11925);
  and g22701 (n11926, n468, n_11416);
  not g22702 (n_11417, n11926);
  and g22703 (n11927, n472, n_11417);
  not g22704 (n_11418, n11927);
  and g22705 (n11928, n476, n_11418);
  not g22706 (n_11419, n11928);
  and g22707 (n11929, n480, n_11419);
  not g22708 (n_11420, n11929);
  and g22709 (n11930, n484, n_11420);
  not g22710 (n_11421, n11930);
  and g22711 (n11931, n488, n_11421);
  not g22712 (n_11422, n11931);
  and g22713 (n11932, n492, n_11422);
  not g22714 (n_11423, n11932);
  and g22715 (n11933, n496, n_11423);
  not g22716 (n_11424, n11933);
  and g22717 (n11934, n500, n_11424);
  not g22718 (n_11425, n11934);
  and g22719 (n11935, n504, n_11425);
  not g22720 (n_11426, n11935);
  and g22721 (n11936, n508, n_11426);
  not g22722 (n_11427, n11936);
  and g22723 (n11937, n512, n_11427);
  not g22724 (n_11428, n11937);
  and g22725 (n11938, n516, n_11428);
  not g22726 (n_11429, n11938);
  and g22727 (n11939, n520, n_11429);
  not g22728 (n_11430, n11939);
  and g22729 (n11940, n524, n_11430);
  not g22730 (n_11431, n11940);
  and g22731 (n11941, n528, n_11431);
  not g22732 (n_11432, n11941);
  and g22733 (n11942, n532, n_11432);
  not g22734 (n_11433, n11942);
  and g22735 (n11943, n536, n_11433);
  not g22736 (n_11434, n11943);
  and g22737 (n11944, n540, n_11434);
  not g22738 (n_11435, n11944);
  and g22739 (n11945, n544, n_11435);
  not g22740 (n_11436, n11945);
  and g22741 (n11946, n548, n_11436);
  not g22742 (n_11437, n11946);
  and g22743 (n11947, n552, n_11437);
  not g22744 (n_11438, n11947);
  and g22745 (n11948, n556, n_11438);
  not g22746 (n_11439, n11948);
  and g22747 (n11949, n560, n_11439);
  not g22748 (n_11440, n11949);
  and g22749 (n11950, n564, n_11440);
  not g22750 (n_11441, n11950);
  and g22751 (n11951, n568, n_11441);
  not g22752 (n_11442, n11951);
  and g22753 (n11952, n572, n_11442);
  not g22754 (n_11443, n11952);
  and g22755 (n11953, n576, n_11443);
  not g22756 (n_11444, n11953);
  and g22757 (n11954, n580, n_11444);
  not g22758 (n_11445, n11954);
  and g22759 (n11955, n584, n_11445);
  not g22760 (n_11446, n11955);
  and g22761 (n11956, n588, n_11446);
  not g22762 (n_11447, n11956);
  and g22763 (n11957, n592, n_11447);
  not g22764 (n_11448, n11957);
  and g22765 (n11958, n596, n_11448);
  not g22766 (n_11449, n11958);
  and g22767 (n11959, n600, n_11449);
  not g22768 (n_11450, n11959);
  and g22769 (n11960, n604, n_11450);
  not g22770 (n_11451, n11960);
  and g22771 (n11961, n608, n_11451);
  not g22772 (n_11452, n11961);
  and g22773 (n11962, n612, n_11452);
  not g22774 (n_11453, n11962);
  and g22775 (n11963, n616, n_11453);
  not g22776 (n_11454, n11963);
  and g22777 (n11964, n620, n_11454);
  not g22778 (n_11455, n11964);
  and g22779 (n11965, n624, n_11455);
  not g22780 (n_11456, n11965);
  and g22781 (n11966, n628, n_11456);
  not g22782 (n_11457, n11966);
  and g22783 (n11967, n632, n_11457);
  not g22784 (n_11458, n11967);
  and g22785 (n11968, n636, n_11458);
  not g22786 (n_11459, n11968);
  and g22787 (n11969, n640, n_11459);
  not g22788 (n_11460, n11969);
  and g22789 (n11970, n644, n_11460);
  not g22790 (n_11461, n11970);
  and g22791 (n11971, n648, n_11461);
  not g22792 (n_11462, n11971);
  and g22793 (n11972, n652, n_11462);
  not g22794 (n_11463, n11972);
  and g22795 (n11973, n656, n_11463);
  not g22796 (n_11464, n11973);
  and g22797 (n11974, n660, n_11464);
  not g22798 (n_11465, n11974);
  and g22799 (n11975, n664, n_11465);
  not g22800 (n_11466, n11975);
  and g22801 (n11976, n668, n_11466);
  not g22802 (n_11467, n11976);
  and g22803 (n11977, n672, n_11467);
  not g22804 (n_11468, n11977);
  and g22805 (n11978, n676, n_11468);
  not g22806 (n_11469, n11978);
  and g22807 (n11979, n680, n_11469);
  not g22808 (n_11470, n11979);
  and g22809 (n11980, n684, n_11470);
  not g22810 (n_11471, n11980);
  and g22811 (n11981, n688, n_11471);
  not g22812 (n_11472, n11981);
  and g22813 (n11982, n692, n_11472);
  not g22814 (n_11473, n11982);
  and g22815 (n11983, n696, n_11473);
  not g22816 (n_11474, n11983);
  and g22817 (n11984, n700, n_11474);
  not g22818 (n_11475, n11984);
  and g22819 (n11985, n704, n_11475);
  not g22820 (n_11476, n11985);
  and g22821 (n11986, n708, n_11476);
  not g22822 (n_11477, n11986);
  and g22823 (n11987, n712, n_11477);
  and g22824 (n11988, \req[125] , n_584);
  not g22825 (n_11478, n11987);
  and g22826 (\grant[125] , n_11478, n11988);
  not g22827 (n_11479, n1058);
  and g22828 (n11990, n_11479, n1483);
  not g22829 (n_11480, n11990);
  and g22830 (n11991, n1486, n_11480);
  not g22831 (n_11481, n11991);
  and g22832 (n11992, n1750, n_11481);
  not g22833 (n_11482, n11992);
  and g22834 (n11993, n731, n_11482);
  not g22835 (n_11483, n11993);
  and g22836 (n11994, n735, n_11483);
  not g22837 (n_11484, n11994);
  and g22838 (n11995, n739, n_11484);
  not g22839 (n_11485, n11995);
  and g22840 (n11996, n743, n_11485);
  not g22841 (n_11486, n11996);
  and g22842 (n11997, n747, n_11486);
  not g22843 (n_11487, n11997);
  and g22844 (n11998, n751, n_11487);
  not g22845 (n_11488, n11998);
  and g22846 (n11999, n755, n_11488);
  not g22847 (n_11489, n11999);
  and g22848 (n12000, n759, n_11489);
  not g22849 (n_11490, n12000);
  and g22850 (n12001, n763, n_11490);
  not g22851 (n_11491, n12001);
  and g22852 (n12002, n767, n_11491);
  not g22853 (n_11492, n12002);
  and g22854 (n12003, n771, n_11492);
  not g22855 (n_11493, n12003);
  and g22856 (n12004, n775, n_11493);
  not g22857 (n_11494, n12004);
  and g22858 (n12005, n779, n_11494);
  not g22859 (n_11495, n12005);
  and g22860 (n12006, n783, n_11495);
  not g22861 (n_11496, n12006);
  and g22862 (n12007, n787, n_11496);
  not g22863 (n_11497, n12007);
  and g22864 (n12008, n791, n_11497);
  not g22865 (n_11498, n12008);
  and g22866 (n12009, n795, n_11498);
  not g22867 (n_11499, n12009);
  and g22868 (n12010, n799, n_11499);
  not g22869 (n_11500, n12010);
  and g22870 (n12011, n803, n_11500);
  not g22871 (n_11501, n12011);
  and g22872 (n12012, n807, n_11501);
  not g22873 (n_11502, n12012);
  and g22874 (n12013, n811, n_11502);
  not g22875 (n_11503, n12013);
  and g22876 (n12014, n815, n_11503);
  not g22877 (n_11504, n12014);
  and g22878 (n12015, n819, n_11504);
  not g22879 (n_11505, n12015);
  and g22880 (n12016, n823, n_11505);
  not g22881 (n_11506, n12016);
  and g22882 (n12017, n827, n_11506);
  not g22883 (n_11507, n12017);
  and g22884 (n12018, n831, n_11507);
  not g22885 (n_11508, n12018);
  and g22886 (n12019, n835, n_11508);
  not g22887 (n_11509, n12019);
  and g22888 (n12020, n839, n_11509);
  not g22889 (n_11510, n12020);
  and g22890 (n12021, n843, n_11510);
  not g22891 (n_11511, n12021);
  and g22892 (n12022, n847, n_11511);
  not g22893 (n_11512, n12022);
  and g22894 (n12023, n851, n_11512);
  not g22895 (n_11513, n12023);
  and g22896 (n12024, n855, n_11513);
  not g22897 (n_11514, n12024);
  and g22898 (n12025, n859, n_11514);
  not g22899 (n_11515, n12025);
  and g22900 (n12026, n863, n_11515);
  not g22901 (n_11516, n12026);
  and g22902 (n12027, n867, n_11516);
  not g22903 (n_11517, n12027);
  and g22904 (n12028, n871, n_11517);
  not g22905 (n_11518, n12028);
  and g22906 (n12029, n875, n_11518);
  not g22907 (n_11519, n12029);
  and g22908 (n12030, n879, n_11519);
  not g22909 (n_11520, n12030);
  and g22910 (n12031, n883, n_11520);
  not g22911 (n_11521, n12031);
  and g22912 (n12032, n887, n_11521);
  not g22913 (n_11522, n12032);
  and g22914 (n12033, n891, n_11522);
  not g22915 (n_11523, n12033);
  and g22916 (n12034, n895, n_11523);
  not g22917 (n_11524, n12034);
  and g22918 (n12035, n899, n_11524);
  not g22919 (n_11525, n12035);
  and g22920 (n12036, n903, n_11525);
  not g22921 (n_11526, n12036);
  and g22922 (n12037, n907, n_11526);
  not g22923 (n_11527, n12037);
  and g22924 (n12038, n911, n_11527);
  not g22925 (n_11528, n12038);
  and g22926 (n12039, n915, n_11528);
  not g22927 (n_11529, n12039);
  and g22928 (n12040, n919, n_11529);
  not g22929 (n_11530, n12040);
  and g22930 (n12041, n923, n_11530);
  not g22931 (n_11531, n12041);
  and g22932 (n12042, n927, n_11531);
  not g22933 (n_11532, n12042);
  and g22934 (n12043, n931, n_11532);
  not g22935 (n_11533, n12043);
  and g22936 (n12044, n935, n_11533);
  not g22937 (n_11534, n12044);
  and g22938 (n12045, n939, n_11534);
  not g22939 (n_11535, n12045);
  and g22940 (n12046, n943, n_11535);
  not g22941 (n_11536, n12046);
  and g22942 (n12047, n947, n_11536);
  not g22943 (n_11537, n12047);
  and g22944 (n12048, n951, n_11537);
  not g22945 (n_11538, n12048);
  and g22946 (n12049, n955, n_11538);
  not g22947 (n_11539, n12049);
  and g22948 (n12050, n959, n_11539);
  not g22949 (n_11540, n12050);
  and g22950 (n12051, n963, n_11540);
  not g22951 (n_11541, n12051);
  and g22952 (n12052, n967, n_11541);
  not g22953 (n_11542, n12052);
  and g22954 (n12053, n971, n_11542);
  not g22955 (n_11543, n12053);
  and g22956 (n12054, n975, n_11543);
  not g22957 (n_11544, n12054);
  and g22958 (n12055, n979, n_11544);
  not g22959 (n_11545, n12055);
  and g22960 (n12056, n983, n_11545);
  not g22961 (n_11546, n12056);
  and g22962 (n12057, n987, n_11546);
  not g22963 (n_11547, n12057);
  and g22964 (n12058, n991, n_11547);
  not g22965 (n_11548, n12058);
  and g22966 (n12059, n995, n_11548);
  not g22967 (n_11549, n12059);
  and g22968 (n12060, n999, n_11549);
  not g22969 (n_11550, n12060);
  and g22970 (n12061, n1003, n_11550);
  not g22971 (n_11551, n12061);
  and g22972 (n12062, n1007, n_11551);
  not g22973 (n_11552, n12062);
  and g22974 (n12063, n1011, n_11552);
  not g22975 (n_11553, n12063);
  and g22976 (n12064, n1015, n_11553);
  not g22977 (n_11554, n12064);
  and g22978 (n12065, n1019, n_11554);
  not g22979 (n_11555, n12065);
  and g22980 (n12066, n1023, n_11555);
  not g22981 (n_11556, n12066);
  and g22982 (n12067, n1027, n_11556);
  not g22983 (n_11557, n12067);
  and g22984 (n12068, n1031, n_11557);
  not g22985 (n_11558, n12068);
  and g22986 (n12069, n1035, n_11558);
  not g22987 (n_11559, n12069);
  and g22988 (n12070, n1039, n_11559);
  not g22989 (n_11560, n12070);
  and g22990 (n12071, n1043, n_11560);
  not g22991 (n_11561, n12071);
  and g22992 (n12072, n1047, n_11561);
  not g22993 (n_11562, n12072);
  and g22994 (n12073, n1051, n_11562);
  and g22995 (n12074, \req[126] , n_845);
  not g22996 (n_11563, n12073);
  and g22997 (\grant[126] , n_11563, n12074);
  not g22998 (n_11564, n1395);
  and g22999 (n12076, n_11564, n1573);
  not g23000 (n_11565, n12076);
  and g23001 (n12077, n1576, n_11565);
  not g23002 (n_11566, n12077);
  and g23003 (n12078, n1837, n_11566);
  not g23004 (n_11567, n12078);
  and g23005 (n12079, n1068, n_11567);
  not g23006 (n_11568, n12079);
  and g23007 (n12080, n1072, n_11568);
  not g23008 (n_11569, n12080);
  and g23009 (n12081, n1076, n_11569);
  not g23010 (n_11570, n12081);
  and g23011 (n12082, n1080, n_11570);
  not g23012 (n_11571, n12082);
  and g23013 (n12083, n1084, n_11571);
  not g23014 (n_11572, n12083);
  and g23015 (n12084, n1088, n_11572);
  not g23016 (n_11573, n12084);
  and g23017 (n12085, n1092, n_11573);
  not g23018 (n_11574, n12085);
  and g23019 (n12086, n1096, n_11574);
  not g23020 (n_11575, n12086);
  and g23021 (n12087, n1100, n_11575);
  not g23022 (n_11576, n12087);
  and g23023 (n12088, n1104, n_11576);
  not g23024 (n_11577, n12088);
  and g23025 (n12089, n1108, n_11577);
  not g23026 (n_11578, n12089);
  and g23027 (n12090, n1112, n_11578);
  not g23028 (n_11579, n12090);
  and g23029 (n12091, n1116, n_11579);
  not g23030 (n_11580, n12091);
  and g23031 (n12092, n1120, n_11580);
  not g23032 (n_11581, n12092);
  and g23033 (n12093, n1124, n_11581);
  not g23034 (n_11582, n12093);
  and g23035 (n12094, n1128, n_11582);
  not g23036 (n_11583, n12094);
  and g23037 (n12095, n1132, n_11583);
  not g23038 (n_11584, n12095);
  and g23039 (n12096, n1136, n_11584);
  not g23040 (n_11585, n12096);
  and g23041 (n12097, n1140, n_11585);
  not g23042 (n_11586, n12097);
  and g23043 (n12098, n1144, n_11586);
  not g23044 (n_11587, n12098);
  and g23045 (n12099, n1148, n_11587);
  not g23046 (n_11588, n12099);
  and g23047 (n12100, n1152, n_11588);
  not g23048 (n_11589, n12100);
  and g23049 (n12101, n1156, n_11589);
  not g23050 (n_11590, n12101);
  and g23051 (n12102, n1160, n_11590);
  not g23052 (n_11591, n12102);
  and g23053 (n12103, n1164, n_11591);
  not g23054 (n_11592, n12103);
  and g23055 (n12104, n1168, n_11592);
  not g23056 (n_11593, n12104);
  and g23057 (n12105, n1172, n_11593);
  not g23058 (n_11594, n12105);
  and g23059 (n12106, n1176, n_11594);
  not g23060 (n_11595, n12106);
  and g23061 (n12107, n1180, n_11595);
  not g23062 (n_11596, n12107);
  and g23063 (n12108, n1184, n_11596);
  not g23064 (n_11597, n12108);
  and g23065 (n12109, n1188, n_11597);
  not g23066 (n_11598, n12109);
  and g23067 (n12110, n1192, n_11598);
  not g23068 (n_11599, n12110);
  and g23069 (n12111, n1196, n_11599);
  not g23070 (n_11600, n12111);
  and g23071 (n12112, n1200, n_11600);
  not g23072 (n_11601, n12112);
  and g23073 (n12113, n1204, n_11601);
  not g23074 (n_11602, n12113);
  and g23075 (n12114, n1208, n_11602);
  not g23076 (n_11603, n12114);
  and g23077 (n12115, n1212, n_11603);
  not g23078 (n_11604, n12115);
  and g23079 (n12116, n1216, n_11604);
  not g23080 (n_11605, n12116);
  and g23081 (n12117, n1220, n_11605);
  not g23082 (n_11606, n12117);
  and g23083 (n12118, n1224, n_11606);
  not g23084 (n_11607, n12118);
  and g23085 (n12119, n1228, n_11607);
  not g23086 (n_11608, n12119);
  and g23087 (n12120, n1232, n_11608);
  not g23088 (n_11609, n12120);
  and g23089 (n12121, n1236, n_11609);
  not g23090 (n_11610, n12121);
  and g23091 (n12122, n1240, n_11610);
  not g23092 (n_11611, n12122);
  and g23093 (n12123, n1244, n_11611);
  not g23094 (n_11612, n12123);
  and g23095 (n12124, n1248, n_11612);
  not g23096 (n_11613, n12124);
  and g23097 (n12125, n1252, n_11613);
  not g23098 (n_11614, n12125);
  and g23099 (n12126, n1256, n_11614);
  not g23100 (n_11615, n12126);
  and g23101 (n12127, n1260, n_11615);
  not g23102 (n_11616, n12127);
  and g23103 (n12128, n1264, n_11616);
  not g23104 (n_11617, n12128);
  and g23105 (n12129, n1268, n_11617);
  not g23106 (n_11618, n12129);
  and g23107 (n12130, n1272, n_11618);
  not g23108 (n_11619, n12130);
  and g23109 (n12131, n1276, n_11619);
  not g23110 (n_11620, n12131);
  and g23111 (n12132, n1280, n_11620);
  not g23112 (n_11621, n12132);
  and g23113 (n12133, n1284, n_11621);
  not g23114 (n_11622, n12133);
  and g23115 (n12134, n1288, n_11622);
  not g23116 (n_11623, n12134);
  and g23117 (n12135, n1292, n_11623);
  not g23118 (n_11624, n12135);
  and g23119 (n12136, n1296, n_11624);
  not g23120 (n_11625, n12136);
  and g23121 (n12137, n1300, n_11625);
  not g23122 (n_11626, n12137);
  and g23123 (n12138, n1304, n_11626);
  not g23124 (n_11627, n12138);
  and g23125 (n12139, n1308, n_11627);
  not g23126 (n_11628, n12139);
  and g23127 (n12140, n1312, n_11628);
  not g23128 (n_11629, n12140);
  and g23129 (n12141, n1316, n_11629);
  not g23130 (n_11630, n12141);
  and g23131 (n12142, n1320, n_11630);
  not g23132 (n_11631, n12142);
  and g23133 (n12143, n1324, n_11631);
  not g23134 (n_11632, n12143);
  and g23135 (n12144, n1328, n_11632);
  not g23136 (n_11633, n12144);
  and g23137 (n12145, n1332, n_11633);
  not g23138 (n_11634, n12145);
  and g23139 (n12146, n1336, n_11634);
  not g23140 (n_11635, n12146);
  and g23141 (n12147, n1340, n_11635);
  not g23142 (n_11636, n12147);
  and g23143 (n12148, n1344, n_11636);
  not g23144 (n_11637, n12148);
  and g23145 (n12149, n1348, n_11637);
  not g23146 (n_11638, n12149);
  and g23147 (n12150, n1352, n_11638);
  not g23148 (n_11639, n12150);
  and g23149 (n12151, n1356, n_11639);
  not g23150 (n_11640, n12151);
  and g23151 (n12152, n1360, n_11640);
  not g23152 (n_11641, n12152);
  and g23153 (n12153, n1364, n_11641);
  not g23154 (n_11642, n12153);
  and g23155 (n12154, n1368, n_11642);
  not g23156 (n_11643, n12154);
  and g23157 (n12155, n1372, n_11643);
  not g23158 (n_11644, n12155);
  and g23159 (n12156, n1376, n_11644);
  not g23160 (n_11645, n12156);
  and g23161 (n12157, n1380, n_11645);
  not g23162 (n_11646, n12157);
  and g23163 (n12158, n1384, n_11646);
  not g23164 (n_11647, n12158);
  and g23165 (n12159, n1388, n_11647);
  and g23166 (n12160, \req[127] , n_1016);
  not g23167 (n_11648, n12159);
  and g23168 (\grant[127] , n_11648, n12160);
  nand g23234 (n_11780, n707, n734, n750, n766);
  nand g23235 (n_11781, n643, n659, n675, n691);
  nand g23236 (n_11782, n846, n862, n878, n894);
  nand g23237 (n_11783, n782, n798, n814, n830);
  nand g23238 (n_11784, n451, n467, n483, n499);
  nand g23239 (n_11785, n388, n403, n419, n435);
  nand g23240 (n_11786, n579, n595, n611, n627);
  nand g23241 (n_11787, n515, n531, n547, n563);
  nand g23242 (n_11788, n1223, n1239, n1255, n1271);
  nand g23243 (n_11789, n1159, n1175, n1191, n1207);
  nand g23244 (n_11790, n1351, n1367, n1383, n1483);
  nand g23245 (n_11791, n1287, n1303, n1319, n1335);
  nand g23246 (n_11792, n974, n990, n1006, n1022);
  nand g23247 (n_11793, n910, n926, n942, n958);
  nand g23248 (n_11794, n1095, n1111, n1127, n1143);
  nand g23249 (n_11795, n1038, n1054, n1064, n1079);
  or g23250 (n_11796, n_11780, n_11781, n_11782, n_11783);
  or g23251 (n_11797, n_11784, n_11785, n_11786, n_11787);
  or g23252 (n_11798, n_11788, n_11789, n_11790, n_11791);
  or g23253 (n_11799, n_11792, n_11793, n_11794, n_11795);
  or g23254 (anyGrant, n_11796, n_11797, n_11798, n_11799);
endmodule

