
module c7552(N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38,
     N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61,
     N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78,
     N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97,
     N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118,
     N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147,
     N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
     N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
     N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
     N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
     N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
     N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
     N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
     N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
     N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263,
     N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299,
     N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334,
     N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367,
     N382, N241_I, N387, N388, N478, N482, N484, N486, N489, N492,
     N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537,
     N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561,
     N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881,
     N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113,
     N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103,
     N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352,
     N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704,
     N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717,
     N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827,
     N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871,
     N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342,
     N241_O);
  input N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41,
       N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
       N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79,
       N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97,
       N100, N103, N106, N109, N110, N111, N112, N113, N114, N115,
       N118, N121, N124, N127, N130, N133, N134, N135, N138, N141,
       N144, N147, N150, N151, N152, N153, N154, N155, N156, N157,
       N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
       N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
       N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
       N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
       N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
       N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
       N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
       N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
       N238, N239, N240, N242, N245, N248, N251, N254, N257, N260,
       N263, N267, N271, N274, N277, N280, N283, N286, N289, N293,
       N296, N299, N303, N307, N310, N313, N316, N319, N322, N325,
       N328, N331, N334, N337, N340, N343, N346, N349, N352, N355,
       N358, N361, N364, N367, N382, N241_I;
  output N387, N388, N478, N482, N484, N486, N489, N492, N501, N505,
       N507, N509, N511, N513, N515, N517, N519, N535, N537, N539,
       N541, N543, N545, N547, N549, N551, N553, N556, N559, N561,
       N563, N565, N567, N569, N571, N573, N582, N643, N707, N813,
       N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112,
       N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102,
       N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351,
       N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641,
       N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716,
       N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763,
       N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870,
       N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340,
       N11342, N241_O;
  wire N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41,
       N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
       N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79,
       N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97,
       N100, N103, N106, N109, N110, N111, N112, N113, N114, N115,
       N118, N121, N124, N127, N130, N133, N134, N135, N138, N141,
       N144, N147, N150, N151, N152, N153, N154, N155, N156, N157,
       N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
       N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
       N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
       N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
       N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
       N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
       N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
       N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
       N238, N239, N240, N242, N245, N248, N251, N254, N257, N260,
       N263, N267, N271, N274, N277, N280, N283, N286, N289, N293,
       N296, N299, N303, N307, N310, N313, N316, N319, N322, N325,
       N328, N331, N334, N337, N340, N343, N346, N349, N352, N355,
       N358, N361, N364, N367, N382, N241_I;
  wire N387, N388, N478, N482, N484, N486, N489, N492, N501, N505,
       N507, N509, N511, N513, N515, N517, N519, N535, N537, N539,
       N541, N543, N545, N547, N549, N551, N553, N556, N559, N561,
       N563, N565, N567, N569, N571, N573, N582, N643, N707, N813,
       N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112,
       N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102,
       N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351,
       N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641,
       N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716,
       N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763,
       N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870,
       N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340,
       N11342, N241_O;
  wire N467, N469, N494, N528, N575, N578, N585, N599;
  wire N604, N609, N628, N641, N642, N644, N651, N660;
  wire N666, N672, N673, N674, N688, N695, N700, N705;
  wire N706, N708, N715, N721, N727, N734, N742, N758;
  wire N759, N762, N768, N774, N780, N786, N794, N800;
  wire N806, N812, N814, N821, N827, N833, N839, N845;
  wire N853, N859, N865, N886, N887, N957, N1028, N1029;
  wire N1109, N1115, N1167, N1222, N1537, N1649, N1708, N1782;
  wire N1793, N1794, N1795, N1796, N1797, N1798, N1811, N1812;
  wire N1813, N1814, N1815, N1816, N1817, N1818, N1819, N1820;
  wire N1821, N1822, N1857, N1858, N1859, N1860, N1861, N1862;
  wire N1863, N1864, N1865, N1866, N1926, N1927, N1928, N1929;
  wire N1930, N1957, N1958, N1959, N1960, N1961, N1962, N1963;
  wire N1966, N1989, N1990, N1991, N1992, N1993, N1994, N1995;
  wire N1996, N2010, N2011, N2012, N2013, N2014, N2064, N2065;
  wire N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073;
  wire N2107, N2108, N2111, N2117, N2171, N2172, N2239, N2241;
  wire N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249;
  wire N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257;
  wire N2268, N2277, N2278, N2279, N2280, N2281, N2299, N2300;
  wire N2301, N2302, N2303, N2321, N2322, N2323, N2324, N2325;
  wire N2337, N2338, N2339, N2340, N2341, N2348, N2349, N2350;
  wire N2351, N2352, N2353, N2354, N2355, N2357, N2358, N2359;
  wire N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367;
  wire N2374, N2375, N2376, N2377, N2378, N2396, N2397, N2398;
  wire N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2418;
  wire N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427;
  wire N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435;
  wire N2436, N2437, N2441, N2446, N2450, N2454, N2458, N2462;
  wire N2466, N2470, N2474, N2478, N2482, N2488, N2496, N2502;
  wire N2508, N2523, N2537, N2538, N2542, N2546, N2550, N2554;
  wire N2561, N2567, N2573, N2604, N2607, N2611, N2615, N2619;
  wire N2626, N2632, N2638, N2644, N2650, N2653, N2654, N2658;
  wire N2662, N2666, N2670, N2674, N2680, N2688, N2692, N2696;
  wire N2700, N2704, N2729, N2733, N2737, N2741, N2745, N2749;
  wire N2753, N2757, N2761, N2766, N2769, N2772, N2775, N2778;
  wire N2781, N2784, N2787, N2790, N2793, N2796, N2866, N2913;
  wire N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921;
  wire N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929;
  wire N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937;
  wire N2988, N3005, N3006, N3007, N3008, N3009, N3020, N3021;
  wire N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029;
  wire N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039;
  wire N3040, N3041, N3073, N3080, N3096, N3097, N3101, N3107;
  wire N3114, N3122, N3126, N3135, N3167, N3168, N3169, N3173;
  wire N3178, N3184, N3185, N3189, N3195, N3202, N3247, N3251;
  wire N3255, N3259, N3263, N3267, N3273, N3281, N3287, N3293;
  wire N3299, N3303, N3307, N3311, N3315, N3322, N3328, N3334;
  wire N3340, N3343, N3349, N3355, N3361, N3362, N3364, N3365;
  wire N3366, N3368, N3370, N3371, N3373, N3375, N3379, N3380;
  wire N3381, N3384, N3390, N3398, N3404, N3410, N3416, N3420;
  wire N3424, N3428, N3432, N3436, N3440, N3444, N3448, N3452;
  wire N3453, N3454, N3458, N3462, N3466, N3470, N3474, N3478;
  wire N3482, N3486, N3507, N3515, N3551, N3552, N3569, N3570;
  wire N3625, N3628, N3781, N3782, N3783, N3786, N3789, N3885;
  wire N3888, N3891, N3953, N3954, N3955, N4193, N4303, N4326;
  wire N4327, N4333, N4334, N4411, N4412, N4463, N4464, N4465;
  wire N4466, N4467, N4468, N4469, N4470, N4471, N4472, N4473;
  wire N4487, N4488, N4490, N4496, N4497, N4498, N4499, N4500;
  wire N4501, N4502, N4503, N4504, N4505, N4506, N4507, N4508;
  wire N4509, N4510, N4511, N4512, N4513, N4515, N4517, N4519;
  wire N4521, N4522, N4523, N4543, N4544, N4545, N4549, N4555;
  wire N4562, N4563, N4566, N4570, N4575, N4611, N4612, N4613;
  wire N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621;
  wire N4622, N4623, N4624, N4625, N4626, N4627, N4628, N4629;
  wire N4630, N4631, N4632, N4633, N4635, N4636, N4637, N4638;
  wire N4640, N4642, N4643, N4645, N4647, N4649, N4651, N4653;
  wire N4656, N4657, N4661, N4667, N4674, N4675, N4678, N4682;
  wire N4687, N4694, N4699, N4700, N4743, N4745, N4746, N4747;
  wire N4748, N4749, N4751, N4756, N4757, N4759, N4760, N4762;
  wire N4766, N4768, N4769, N4776, N4781, N4782, N4783, N4784;
  wire N4795, N4803, N4806, N4813, N4844, N4940, N4997, N5030;
  wire N5165, N5167, N5168, N5169, N5170, N5171, N5177, N5178;
  wire N5179, N5180, N5181, N5182, N5183, N5184, N5185, N5186;
  wire N5187, N5188, N5189, N5190, N5191, N5192, N5193, N5196;
  wire N5197, N5198, N5199, N5200, N5201, N5202, N5203, N5204;
  wire N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290;
  wire N5291, N5292, N5293, N5294, N5295, N5296, N5297, N5298;
  wire N5299, N5300, N5314, N5315, N5316, N5317, N5318, N5319;
  wire N5320, N5321, N5322, N5323, N5324, N5363, N5364, N5365;
  wire N5366, N5367, N5425, N5426, N5427, N5429, N5430, N5431;
  wire N5432, N5433, N5451, N5452, N5453, N5454, N5455, N5456;
  wire N5457, N5469, N5474, N5475, N5476, N5477, N5571, N5572;
  wire N5573, N5574, N5584, N5585, N5586, N5587, N5602, N5603;
  wire N5604, N5605, N5631, N5632, N5640, N5654, N5670, N5683;
  wire N5735, N5736, N5740, N5744, N5747, N5751, N5755, N5758;
  wire N5762, N5766, N5769, N5770, N5771, N5778, N5789, N5799;
  wire N5807, N5821, N5837, N5850, N5856, N5943, N5944, N5945;
  wire N5946, N5947, N5948, N5949, N5950, N5951, N5952, N5953;
  wire N5954, N5955, N5956, N5957, N5958, N5959, N5960, N5966;
  wire N5991, N5996, N6000, N6003, N6009, N6014, N6018, N6021;
  wire N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029;
  wire N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037;
  wire N6038, N6039, N6040, N6041, N6047, N6052, N6056, N6059;
  wire N6060, N6061, N6062, N6063, N6064, N6065, N6066, N6067;
  wire N6068, N6069, N6070, N6071, N6072, N6073, N6074, N6075;
  wire N6076, N6077, N6078, N6079, N6083, N6087, N6091, N6096;
  wire N6097, N6102, N6122, N6125, N6127, N6131, N6135, N6136;
  wire N6137, N6141, N6145, N6148, N6149, N6150, N6151, N6152;
  wire N6153, N6154, N6156, N6157, N6158, N6159, N6160, N6161;
  wire N6162, N6163, N6164, N6165, N6166, N6170, N6174, N6177;
  wire N6186, N6191, N6192, N6194, N6195, N6196, N6199, N6203;
  wire N6217, N6235, N6243, N6246, N6249, N6252, N6263, N6266;
  wire N6540, N6541, N6542, N6543, N6544, N6545, N6546, N6547;
  wire N6594, N6595, N6596, N6597, N6598, N6599, N6600, N6601;
  wire N6602, N6603, N6604, N6605, N6606, N6621, N6622, N6623;
  wire N6624, N6625, N6626, N6627, N6628, N6629, N6639, N6640;
  wire N6641, N6642, N6643, N6644, N6645, N6646, N6647, N6648;
  wire N6658, N6659, N6660, N6661, N6668, N6677, N6678, N6679;
  wire N6680, N6681, N6682, N6683, N6684, N6685, N6686, N6687;
  wire N6688, N6689, N6690, N6702, N6703, N6704, N6705, N6706;
  wire N6707, N6708, N6709, N6710, N6711, N6712, N6729, N6730;
  wire N6731, N6732, N6733, N6734, N6735, N6736, N6741, N6742;
  wire N6743, N6744, N6751, N6752, N6753, N6754, N6755, N6756;
  wire N6757, N6758, N6761, N6762, N6766, N6767, N6768, N6769;
  wire N6770, N6771, N6772, N6773, N6777, N6778, N6779, N6782;
  wire N6783, N6784, N6797, N6800, N6803, N6806, N6809, N6812;
  wire N6833, N6836, N6837, N6838, N6839, N6840, N6841, N6844;
  wire N6845, N6848, N6849, N6850, N6851, N6852, N6853, N6854;
  wire N6855, N6859, N6860, N6861, N6864, N6865, N6866, N6881;
  wire N6894, N6901, N6912, N6923, N6929, N6936, N6946, N6957;
  wire N6967, N6968, N6969, N7057, N7060, N7061, N7062, N7064;
  wire N7065, N7066, N7067, N7068, N7073, N7077, N7080, N7086;
  wire N7091, N7095, N7098, N7099, N7100, N7103, N7104, N7105;
  wire N7106, N7107, N7114, N7125, N7136, N7142, N7149, N7159;
  wire N7170, N7180, N7187, N7188, N7191, N7194, N7198, N7202;
  wire N7205, N7209, N7213, N7314, N7318, N7322, N7325, N7328;
  wire N7331, N7334, N7337, N7346, N7351, N7355, N7358, N7364;
  wire N7369, N7373, N7376, N7377, N7378, N7381, N7384, N7387;
  wire N7391, N7394, N7398, N7402, N7441, N7444, N7477, N7478;
  wire N7552, N7556, N7557, N7558, N7559, N7560, N7563, N7566;
  wire N7569, N7573, N7574, N7577, N7580, N7581, N7582, N7585;
  wire N7588, N7591, N7609, N7613, N7649, N7650, N7655, N7659;
  wire N7744, N7825, N7826, N7852, N8114, N8117, N8131, N8134;
  wire N8144, N8145, N8146, N8156, N8166, N8169, N8183, N8186;
  wire N8204, N8208, N8216, N8217, N8218, N8219, N8232, N8233;
  wire N8242, N8243, N8244, N8245, N8246, N8247, N8248, N8249;
  wire N8250, N8251, N8252, N8253, N8254, N8262, N8269, N8274;
  wire N8276, N8278, N8280, N8281, N8282, N8283, N8284, N8285;
  wire N8288, N8294, N8298, N8307, N8315, N8322, N8323, N8324;
  wire N8326, N8333, N8337, N8338, N8339, N8340, N8341, N8342;
  wire N8345, N8346, N8348, N8349, N8350, N8351, N8352, N8353;
  wire N8354, N8355, N8356, N8357, N8394, N8404, N8405, N8409;
  wire N8410, N8411, N8412, N8415, N8416, N8417, N8418, N8421;
  wire N8430, N8433, N8434, N8435, N8436, N8437, N8438, N8441;
  wire N8442, N8444, N8447, N8448, N8449, N8450, N8451, N8452;
  wire N8453, N8454, N8455, N8456, N8457, N8460, N8463, N8466;
  wire N8469, N8483, N8484, N8497, N8507, N8513, N8518, N8519;
  wire N8522, N8537, N8539, N8540, N8541, N8545, N8546, N8547;
  wire N8548, N8551, N8552, N8553, N8554, N8555, N8558, N8561;
  wire N8564, N8578, N8579, N8607, N8608, N8609, N8610, N8627;
  wire N8717, N8727, N8730, N8733, N8734, N8753, N8754, N8755;
  wire N8756, N8811, N8814, N8815, N8816, N8817, N8818, N8857;
  wire N8861, N8862, N8863, N8864, N8865, N8866, N8871, N8874;
  wire N8879, N8880, N8881, N8882, N8883, N8884, N8886, N8887;
  wire N8888, N8898, N8902, N8924, N8931, N8943, N8950, N8956;
  wire N8959, N8960, N8963, N8966, N8991, N8992, N8996, N9005;
  wire N9024, N9025, N9029, N9035, N9053, N9054, N9064, N9065;
  wire N9066, N9067, N9068, N9071, N9072, N9073, N9074, N9077;
  wire N9079, N9087, N9088, N9089, N9092, N9093, N9094, N9095;
  wire N9098, N9099, N9103, N9107, N9111, N9146, N9149, N9159;
  wire N9160, N9161, N9165, N9169, N9173, N9179, N9180, N9181;
  wire N9182, N9203, N9206, N9220, N9223, N9234, N9235, N9236;
  wire N9237, N9243, N9244, N9245, N9246, N9247, N9248, N9249;
  wire N9250, N9251, N9252, N9256, N9257, N9258, N9259, N9260;
  wire N9261, N9262, N9265, N9271, N9272, N9273, N9274, N9275;
  wire N9276, N9280, N9285, N9286, N9287, N9288, N9290, N9294;
  wire N9297, N9298, N9299, N9307, N9314, N9315, N9318, N9323;
  wire N9324, N9326, N9332, N9344, N9352, N9356, N9359, N9360;
  wire N9361, N9363, N9365, N9367, N9368, N9369, N9370, N9371;
  wire N9372, N9375, N9385, N9392, N9394, N9396, N9397, N9398;
  wire N9399, N9400, N9401, N9402, N9407, N9408, N9412, N9413;
  wire N9415, N9417, N9418, N9419, N9420, N9421, N9422, N9426;
  wire N9429, N9432, N9435, N9442, N9445, N9478, N9485, N9488;
  wire N9517, N9520, N9526, N9539, N9540, N9541, N9543, N9551;
  wire N9555, N9556, N9557, N9560, N9561, N9562, N9563, N9564;
  wire N9565, N9566, N9568, N9569, N9570, N9575, N9581, N9582;
  wire N9585, N9591, N9592, N9593, N9594, N9595, N9596, N9597;
  wire N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9608;
  wire N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9621;
  wire N9622, N9623, N9624, N9626, N9629, N9632, N9635, N9642;
  wire N9645, N9646, N9650, N9653, N9656, N9659, N9660, N9662;
  wire N9663, N9666, N9667, N9671, N9679, N9682, N9685, N9690;
  wire N9691, N9692, N9695, N9698, N9702, N9707, N9715, N9716;
  wire N9717, N9720, N9721, N9722, N9723, N9726, N9727, N9732;
  wire N9733, N9734, N9736, N9737, N9738, N9739, N9740, N9741;
  wire N9742, N9754, N9758, N9762, N9763, N9764, N9765, N9766;
  wire N9767, N9768, N9769, N9773, N9775, N9784, N9785, N9786;
  wire N9790, N9791, N9795, N9796, N9797, N9798, N9799, N9800;
  wire N9801, N9802, N9803, N9805, N9806, N9813, N9814, N9815;
  wire N9816, N9817, N9820, N9825, N9826, N9827, N9828, N9829;
  wire N9830, N9835, N9836, N9837, N9838, N9846, N9847, N9863;
  wire N9873, N9876, N9890, N9891, N9892, N9893, N9894, N9895;
  wire N9896, N9897, N9898, N9899, N9900, N9901, N9902, N9903;
  wire N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911;
  wire N9917, N9923, N9924, N9925, N9932, N9935, N9938, N9939;
  wire N9945, N9946, N9947, N9948, N9949, N9953, N9954, N9955;
  wire N9956, N9957, N9958, N9959, N9960, N9961, N9964, N9967;
  wire N9968, N9969, N9970, N9971, N9972, N9974, N9975, N9976;
  wire N9977, N9978, N9979, N9983, N9986, N9989, N9992, N9995;
  wire N9996, N9998, N9999, N10002, N10003, N10007, N10010, N10013;
  wire N10014, N10015, N10016, N10017, N10020, N10021, N10022, N10023;
  wire N10024, N10026, N10028, N10032, N10033, N10034, N10035, N10036;
  wire N10037, N10038, N10039, N10040, N10041, N10042, N10043, N10050;
  wire N10053, N10054, N10055, N10056, N10057, N10058, N10059, N10060;
  wire N10061, N10062, N10067, N10070, N10073, N10076, N10077, N10082;
  wire N10083, N10084, N10085, N10086, N10093, N10094, N10105, N10106;
  wire N10107, N10108, N10113, N10114, N10115, N10116, N10119, N10124;
  wire N10130, N10131, N10132, N10133, N10134, N10135, N10136, N10137;
  wire N10138, N10139, N10140, N10141, N10148, N10155, N10156, N10157;
  wire N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165;
  wire N10170, N10173, N10176, N10177, N10178, N10179, N10180, N10183;
  wire N10186, N10189, N10192, N10195, N10196, N10197, N10200, N10203;
  wire N10204, N10205, N10206, N10212, N10213, N10230, N10231, N10232;
  wire N10233, N10234, N10237, N10238, N10239, N10240, N10241, N10242;
  wire N10247, N10248, N10259, N10264, N10265, N10266, N10267, N10268;
  wire N10269, N10270, N10271, N10272, N10278, N10279, N10280, N10281;
  wire N10282, N10283, N10287, N10288, N10289, N10290, N10291, N10292;
  wire N10293, N10294, N10295, N10296, N10299, N10300, N10301, N10306;
  wire N10307, N10314, N10315, N10316, N10317, N10318, N10321, N10324;
  wire N10325, N10326, N10327, N10328, N10329, N10330, N10331, N10332;
  wire N10333, N10334, N10337, N10338, N10339, N10340, N10341, N10344;
  wire N10354, N10357, N10360, N10367, N10375, N10381, N10388, N10391;
  wire N10399, N10402, N10406, N10409, N10412, N10415, N10419, N10422;
  wire N10425, N10428, N10431, N10432, N10437, N10438, N10439, N10440;
  wire N10441, N10444, N10445, N10450, N10451, N10455, N10456, N10465;
  wire N10466, N10479, N10497, N10509, N10512, N10515, N10516, N10517;
  wire N10518, N10519, N10522, N10525, N10528, N10531, N10534, N10535;
  wire N10536, N10539, N10542, N10543, N10544, N10545, N10546, N10547;
  wire N10548, N10549, N10550, N10551, N10552, N10553, N10554, N10555;
  wire N10556, N10557, N10558, N10559, N10560, N10561, N10562, N10563;
  wire N10564, N10565, N10566, N10567, N10568, N10569, N10570, N10571;
  wire N10572, N10573, N10577, N10581, N10582, N10583, N10587, N10588;
  wire N10589, N10594, N10595, N10596, N10597, N10598, N10609, N10610;
  wire N10621, N10626, N10627, N10629, N10631, N10637, N10638, N10639;
  wire N10640, N10642, N10643, N10644, N10645, N10647, N10648, N10649;
  wire N10652, N10659, N10662, N10665, N10668, N10671, N10672, N10673;
  wire N10674, N10675, N10678, N10681, N10682, N10683, N10684, N10685;
  wire N10686, N10687, N10688, N10689, N10690, N10691, N10694, N10695;
  wire N10696, N10697, N10698, N10701, N10705, N10707, N10708, N10709;
  wire N10710, N10719, N10720, N10730, N10731, N10737, N10738, N10739;
  wire N10746, N10747, N10748, N10749, N10750, N10753, N10754, N10764;
  wire N10765, N10766, N10767, N10768, N10769, N10770, N10771, N10772;
  wire N10773, N10774, N10775, N10776, N10784, N10789, N10792, N10796;
  wire N10797, N10798, N10799, N10800, N10803, N10806, N10809, N10812;
  wire N10815, N10816, N10817, N10820, N10823, N10824, N10825, N10826;
  wire N10832, N10833, N10834, N10835, N10836, N10845, N10846, N10857;
  wire N10862, N10863, N10864, N10865, N10866, N10867, N10872, N10873;
  wire N10874, N10875, N10876, N10879, N10882, N10883, N10884, N10885;
  wire N10886, N10887, N10888, N10889, N10890, N10891, N10892, N10895;
  wire N10896, N10897, N10898, N10899, N10902, N10909, N10910, N10915;
  wire N10916, N10917, N10918, N10919, N10922, N10923, N10928, N10931;
  wire N10934, N10935, N10936, N10937, N10938, N10941, N10944, N10947;
  wire N10950, N10953, N10954, N10955, N10958, N10961, N10962, N10963;
  wire N10964, N10969, N10970, N10981, N10986, N10987, N10988, N10989;
  wire N10990, N10991, N10992, N10995, N10998, N10999, N11000, N11001;
  wire N11002, N11003, N11004, N11005, N11006, N11007, N11008, N11011;
  wire N11012, N11013, N11014, N11015, N11018, N11023, N11024, N11027;
  wire N11028, N11029, N11030, N11031, N11034, N11035, N11040, N11041;
  wire N11042, N11043, N11044, N11047, N11050, N11053, N11056, N11059;
  wire N11062, N11065, N11066, N11067, N11070, N11073, N11074, N11075;
  wire N11076, N11077, N11078, N11095, N11098, N11099, N11100, N11103;
  wire N11106, N11107, N11108, N11109, N11110, N11111, N11112, N11113;
  wire N11114, N11115, N11116, N11117, N11118, N11119, N11120, N11121;
  wire N11122, N11123, N11124, N11127, N11130, N11137, N11138, N11139;
  wire N11140, N11141, N11142, N11143, N11144, N11145, N11152, N11153;
  wire N11154, N11155, N11156, N11159, N11162, N11165, N11168, N11171;
  wire N11174, N11177, N11180, N11183, N11184, N11185, N11186, N11187;
  wire N11188, N11205, N11210, N11211, N11212, N11213, N11214, N11215;
  wire N11216, N11217, N11218, N11219, N11220, N11222, N11223, N11224;
  wire N11225, N11226, N11227, N11228, N11229, N11231, N11232, N11233;
  wire N11236, N11239, N11242, N11243, N11244, N11245, N11246, N11250;
  wire N11252, N11257, N11260, N11261, N11262, N11263, N11264, N11265;
  wire N11267, N11268, N11269, N11270, N11272, N11277, N11278, N11279;
  wire N11280, N11282, N11283, N11284, N11285, N11286, N11288, N11289;
  wire N11290, N11291, N11292, N11293, N11294, N11295, N11296, N11297;
  wire N11298, N11299, N11302, N11307, N11308, N11309, N11312, N11313;
  wire N11314, N11315, N11316, N11317, N11320, N11321, N11323, N11327;
  wire N11328, N11329, N11331, N11335, N11336, N11337, N11338, N11339;
  wire N11341, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_346, n_347;
  wire n_348, n_349, n_350, n_352, n_353, n_358, n_360, n_362;
  wire n_364;
  assign N-241_O = N241_I;
  assign N-10840 = N10839;
  assign N10838 = N10837;
  assign N10103 = N10102;
  assign N1490 = N1;
  assign N1489 = N1113;
  assign N1114 = N582;
  assign N1112 = N1110;
  assign N1111 = N582;
  assign N945 = N106;
  assign N889 = N1;
  assign N813 = N340;
  assign N707 = N277;
  assign N643 = N251;
  assign N573 = N364;
  assign N571 = N361;
  assign N569 = N358;
  assign N567 = N355;
  assign N565 = N352;
  assign N563 = N349;
  assign N561 = N346;
  assign N559 = N343;
  assign N556 = N337;
  assign N553 = N334;
  assign N551 = N331;
  assign N549 = N328;
  assign N547 = N325;
  assign N545 = N322;
  assign N543 = N319;
  assign N541 = N316;
  assign N539 = N313;
  assign N537 = N310;
  assign N535 = N307;
  assign N519 = N303;
  assign N517 = N299;
  assign N515 = N296;
  assign N513 = N293;
  assign N511 = N289;
  assign N509 = N286;
  assign N507 = N283;
  assign N505 = N280;
  assign N501 = N274;
  assign N492 = N267;
  assign N489 = N263;
  assign N486 = N260;
  assign N484 = N257;
  assign N482 = N254;
  assign N478 = N248;
  assign N388 = N1;
  assign N387 = N1;
  and AND2_4 (N469, N134, N133);
  and AND2_69 (N688, N382, N263);
  and AND2_113 (N886, N528, N578);
  and AND2_114 (N887, N575, N494);
  and AND2_118 (N1028, N382, N641);
  and AND2_120 (N1109, N469, N585);
  and AND2_136 (N1167, N700, N38);
  and AND2_226 (N1537, N957, N38);
  and AND2_228 (N1649, N1029, N38);
  and AND2_234 (N1781, N163, N1);
  and AND2_235 (N1782, N170, N18);
  and AND2_238 (N1793, N169, N18);
  and AND2_239 (N1794, N168, N18);
  and AND2_240 (N1795, N167, N18);
  and AND2_241 (N1796, N166, N18);
  and AND2_242 (N1797, N165, N18);
  and AND2_243 (N1798, N164, N18);
  and AND2_246 (N1811, N177, N18);
  and AND2_247 (N1812, N176, N18);
  and AND2_248 (N1813, N175, N18);
  and AND2_249 (N1814, N174, N18);
  and AND2_250 (N1815, N173, N18);
  and AND2_251 (N1816, N157, N18);
  and AND2_252 (N1817, N156, N18);
  and AND2_253 (N1818, N155, N18);
  and AND2_254 (N1819, N154, N18);
  and AND2_255 (N1820, N153, N18);
  and AND2_272 (N1857, N181, N18);
  and AND2_273 (N1858, N171, N18);
  and AND2_274 (N1859, N180, N18);
  and AND2_275 (N1860, N179, N18);
  and AND2_276 (N1861, N178, N18);
  and AND2_277 (N1862, N161, N18);
  and AND2_278 (N1863, N151, N18);
  and AND2_279 (N1864, N160, N18);
  and AND2_280 (N1865, N159, N18);
  and AND2_281 (N1866, N158, N18);
  and AND2_306 (N1926, N44, N695);
  and AND2_307 (N1927, N41, N695);
  and AND2_308 (N1928, N29, N695);
  and AND2_309 (N1929, N26, N695);
  and AND2_310 (N1930, N23, N695);
  and AND2_329 (N1957, N209, N18);
  and AND2_330 (N1958, N216, N18);
  and AND2_331 (N1959, N215, N18);
  and AND2_332 (N1960, N214, N18);
  and AND2_333 (N1961, N213, N18);
  and AND2_334 (N1962, N212, N18);
  and AND2_335 (N1963, N211, N18);
  and AND2_337 (N1966, N1222, N38);
  and AND2_350 (N1989, N642, N18);
  and AND2_351 (N1990, N644, N18);
  and AND2_352 (N1991, N651, N18);
  and AND2_353 (N1992, N674, N18);
  and AND2_354 (N1993, N660, N18);
  and AND2_355 (N1994, N666, N18);
  and AND2_356 (N1995, N672, N18);
  and AND2_357 (N1996, N673, N18);
  and AND2_360 (N2010, N47, N695);
  and AND2_361 (N2011, N35, N695);
  and AND2_362 (N2012, N32, N695);
  and AND2_363 (N2013, N50, N695);
  and AND2_364 (N2014, N66, N695);
  and AND2_380 (N2064, N706, N18);
  and AND2_381 (N2065, N708, N18);
  and AND2_382 (N2066, N715, N18);
  and AND2_383 (N2067, N721, N18);
  and AND2_384 (N2068, N727, N18);
  and AND2_385 (N2069, N599, N18);
  and AND2_386 (N2070, N734, N18);
  and AND2_387 (N2071, N742, N18);
  and AND2_388 (N2072, N604, N18);
  and AND2_389 (N2073, N609, N18);
  and AND2_431 (N2277, N141, N695);
  and AND2_432 (N2278, N147, N695);
  and AND2_433 (N2279, N138, N695);
  and AND2_434 (N2280, N144, N695);
  and AND2_435 (N2281, N135, N695);
  and AND2_443 (N2299, N103, N695);
  and AND2_444 (N2300, N130, N695);
  and AND2_445 (N2301, N127, N695);
  and AND2_446 (N2302, N124, N695);
  and AND2_447 (N2303, N100, N695);
  and AND2_455 (N2321, N115, N695);
  and AND2_456 (N2322, N118, N695);
  and AND2_457 (N2323, N97, N695);
  and AND2_458 (N2324, N94, N695);
  and AND2_459 (N2325, N121, N695);
  and AND2_466 (N2337, N208, N18);
  and AND2_467 (N2338, N198, N18);
  and AND2_468 (N2339, N207, N18);
  and AND2_469 (N2340, N206, N18);
  and AND2_470 (N2341, N205, N18);
  and AND2_487 (N2358, N114, N695);
  and AND2_488 (N2359, N113, N695);
  and AND2_489 (N2360, N111, N695);
  and AND2_490 (N2361, N87, N695);
  and AND2_491 (N2362, N112, N695);
  and AND2_492 (N2363, N88, N695);
  and AND2_493 (N2364, N245, N695);
  and AND2_494 (N2365, N271, N695);
  and AND2_495 (N2366, N759, N695);
  and AND2_496 (N2367, N70, N695);
  and AND2_498 (N2374, N193, N18);
  and AND2_499 (N2375, N192, N18);
  and AND2_500 (N2376, N191, N18);
  and AND2_501 (N2377, N190, N18);
  and AND2_502 (N2378, N189, N18);
  and AND2_510 (N2396, N58, N695);
  and AND2_511 (N2397, N77, N695);
  and AND2_512 (N2398, N78, N695);
  and AND2_513 (N2399, N59, N695);
  and AND2_514 (N2400, N81, N695);
  and AND2_515 (N2401, N80, N695);
  and AND2_516 (N2402, N79, N695);
  and AND2_517 (N2403, N60, N695);
  and AND2_518 (N2404, N61, N695);
  and AND2_519 (N2405, N62, N695);
  and AND2_522 (N2418, N69, N695);
  and AND2_524 (N2420, N74, N695);
  and AND2_525 (N2421, N76, N695);
  and AND2_526 (N2422, N75, N695);
  and AND2_527 (N2423, N73, N695);
  and AND2_528 (N2424, N53, N695);
  and AND2_529 (N2425, N54, N695);
  and AND2_530 (N2426, N55, N695);
  and AND2_531 (N2427, N56, N695);
  and AND2_532 (N2428, N82, N695);
  and AND2_533 (N2429, N65, N695);
  and AND2_534 (N2430, N83, N695);
  and AND2_535 (N2431, N84, N695);
  and AND2_536 (N2432, N85, N695);
  and AND2_537 (N2433, N64, N695);
  and AND2_538 (N2434, N63, N695);
  and AND2_539 (N2435, N86, N695);
  and AND2_540 (N2436, N109, N695);
  and AND2_541 (N2437, N110, N695);
  and AND2_542 (N2441, N2239, N628);
  and AND2_544 (N2446, N2241, N628);
  and AND2_545 (N2450, N2242, N628);
  and AND2_546 (N2454, N2243, N628);
  and AND2_547 (N2458, N2244, N628);
  and AND2_548 (N2462, N2247, N628);
  and AND2_549 (N2466, N2248, N628);
  and AND2_550 (N2470, N2249, N628);
  and AND2_551 (N2474, N2250, N628);
  and AND2_552 (N2478, N2251, N628);
  and AND2_553 (N2482, N2252, N628);
  and AND2_554 (N2488, N2253, N628);
  and AND2_555 (N2496, N2254, N628);
  and AND2_556 (N2502, N2255, N628);
  and AND2_557 (N2508, N2256, N628);
  and AND2_573 (N2619, N2348, N628);
  and AND2_574 (N2626, N2349, N628);
  and AND2_575 (N2632, N2350, N628);
  and AND2_576 (N2638, N2351, N628);
  and AND2_577 (N2644, N2352, N628);
  and AND2_603 (N2766, N2354, N628);
  and AND2_604 (N2769, N2353, N628);
  and AND2_605 (N2772, N2246, N628);
  and AND2_606 (N2775, N2245, N628);
  and AND2_614 (N2866, N2257, N1537);
  and AND2_619 (N2913, N204, N18);
  and AND2_620 (N2914, N203, N18);
  and AND2_621 (N2915, N202, N18);
  and AND2_622 (N2916, N201, N18);
  and AND2_623 (N2917, N200, N18);
  and AND2_624 (N2918, N235, N18);
  and AND2_625 (N2919, N234, N18);
  and AND2_626 (N2920, N233, N18);
  and AND2_627 (N2921, N232, N18);
  and AND2_628 (N2922, N231, N18);
  and AND2_629 (N2923, N197, N18);
  and AND2_630 (N2924, N187, N18);
  and AND2_631 (N2925, N196, N18);
  and AND2_632 (N2926, N195, N18);
  and AND2_633 (N2927, N194, N18);
  and AND2_634 (N2928, N227, N18);
  and AND2_635 (N2929, N217, N18);
  and AND2_636 (N2930, N226, N18);
  and AND2_637 (N2931, N225, N18);
  and AND2_638 (N2932, N224, N18);
  and AND2_639 (N2933, N239, N18);
  and AND2_640 (N2934, N229, N18);
  and AND2_641 (N2935, N238, N18);
  and AND2_642 (N2936, N237, N18);
  and AND2_643 (N2937, N236, N18);
  and AND2_645 (N3005, N223, N18);
  and AND2_646 (N3006, N222, N18);
  and AND2_647 (N3007, N221, N18);
  and AND2_648 (N3008, N220, N18);
  and AND2_649 (N3009, N219, N18);
  and AND2_650 (N3020, N812, N18);
  and AND2_651 (N3021, N814, N18);
  and AND2_652 (N3022, N821, N18);
  and AND2_653 (N3023, N827, N18);
  and AND2_654 (N3024, N833, N18);
  and AND2_655 (N3025, N839, N18);
  and AND2_656 (N3026, N845, N18);
  and AND2_657 (N3027, N853, N18);
  and AND2_658 (N3028, N859, N18);
  and AND2_659 (N3029, N865, N18);
  and AND2_660 (N3032, N758, N18);
  and AND2_661 (N3033, N759, N18);
  and AND2_662 (N3034, N762, N18);
  and AND2_663 (N3035, N768, N18);
  and AND2_664 (N3036, N774, N18);
  and AND2_665 (N3037, N780, N18);
  and AND2_666 (N3038, N786, N18);
  and AND2_667 (N3039, N794, N18);
  and AND2_668 (N3040, N800, N18);
  and AND2_669 (N3041, N806, N18);
  and AND2_676 (N3096, N666, N2644);
  and AND2_677 (N3097, N660, N2638);
  and AND2_678 (N3101, N674, N2632);
  and AND2_679 (N3107, N651, N2626);
  and AND2_680 (N3114, N644, N2619);
  and AND2_681 (N3122, N2523, N2257);
  and AND2_695 (N3168, N609, N2508);
  and AND2_696 (N3169, N604, N2502);
  and AND2_697 (N3173, N742, N2496);
  and AND2_698 (N3178, N734, N2488);
  and AND2_699 (N3184, N599, N2482);
  and AND2_700 (N3185, N727, N2573);
  and AND2_701 (N3189, N721, N2567);
  and AND2_702 (N3195, N715, N2561);
  and AND2_703 (N3202, N708, N2554);
  and AND2_735 (N3361, N2761, N2478);
  and AND2_736 (N3362, N2757, N2474);
  and AND2_738 (N3364, N2749, N2466);
  and AND2_739 (N3365, N2745, N2462);
  and AND2_740 (N3366, N2741, N2550);
  and AND2_742 (N3368, N2733, N2542);
  and AND2_744 (N3370, N2670, N2458);
  and AND2_745 (N3371, N2666, N2454);
  and AND2_747 (N3373, N2658, N2446);
  and AND2_749 (N3375, N2988, N2650);
  and AND2_750 (N3379, N2650, N1966);
  and AND2_752 (N3381, N695, N2604);
  and AND2_1012 (N4544, N806, N3293);
  and AND2_1013 (N4545, N800, N3287);
  and AND2_1014 (N4549, N794, N3281);
  and AND2_1015 (N4555, N3273, N786);
  and AND2_1016 (N4562, N780, N3267);
  and AND2_1017 (N4563, N774, N3355);
  and AND2_1018 (N4566, N768, N3349);
  and AND2_1019 (N4570, N762, N3343);
  and AND2_1049 (N4630, N3448, N2704);
  and AND2_1051 (N4632, N3444, N2700);
  and AND2_1054 (N4635, N3436, N2692);
  and AND2_1056 (N4637, N3432, N2688);
  and AND2_1057 (N4638, N3428, N3311);
  and AND2_1059 (N4640, N3420, N3303);
  and AND2_1073 (N4656, N865, N3410);
  and AND2_1074 (N4657, N859, N3404);
  and AND2_1075 (N4661, N853, N3398);
  and AND2_1076 (N4667, N3390, N845);
  and AND2_1077 (N4674, N839, N3384);
  and AND2_1078 (N4675, N833, N3334);
  and AND2_1079 (N4678, N827, N3328);
  and AND2_1080 (N4682, N821, N3322);
  and AND2_1081 (N4687, N814, N3315);
  and AND2_1112 (N4756, N3482, N3263);
  and AND2_1113 (N4757, N3478, N3259);
  and AND2_1115 (N4759, N3470, N3251);
  and AND2_1116 (N4760, N3466, N3247);
  and AND2_1118 (N4762, N3462, N2615);
  and AND2_1122 (N4766, N3454, N2607);
  and AND2_1125 (N4769, N3340, N695);
  and AND2_1447 (N5960, N2674, N4769);
  and AND2_1751 (N6766, N5632, N3097);
  and AND2_1755 (N6770, N5640, N3101);
  and AND2_1762 (N6777, N5654, N3107);
  and AND2_1767 (N6782, N5670, N3114);
  and AND2_1768 (N6783, N5683, N5670);
  and AND2_1793 (N6836, N5771, N3169);
  and AND2_1796 (N6839, N5778, N3173);
  and AND2_1801 (N6844, N5789, N3178);
  and AND2_1803 (N6848, N5799, N3185);
  and AND2_1807 (N6852, N5807, N3189);
  and AND2_1814 (N6859, N5821, N3195);
  and AND2_1819 (N6864, N5837, N3202);
  and AND2_1820 (N6865, N5850, N5789);
  and AND2_1821 (N6866, N5856, N5837);
  and AND2_1867 (N7060, N5991, N3362);
  and AND2_1871 (N7064, N6003, N3366);
  and AND2_1885 (N7103, N6041, N3371);
  and AND2_2067 (N8262, N3122, N6762);
  and AND2_2068 (N8269, N3122, N6784);
  and AND2_2086 (N8298, N6833, N6845);
  and AND2_2087 (N8307, N6833, N6881);
  and AND2_2098 (N8337, N6894, N4545);
  and AND2_2101 (N8340, N6901, N4549);
  and AND2_2106 (N8345, N6912, N4555);
  and AND2_2107 (N8346, N6923, N6912);
  and AND2_2109 (N8348, N6929, N4563);
  and AND2_2113 (N8352, N6936, N4566);
  and AND2_2116 (N8355, N4570, N6946);
  and AND2_2118 (N8357, N6957, N5960);
  and AND2_2147 (N8404, N7057, N7826);
  and AND2_2149 (N8409, N7068, N4632);
  and AND2_2153 (N8415, N7080, N4638);
  and AND2_2157 (N8421, N3375, N7100);
  and AND2_2159 (N8433, N7107, N4657);
  and AND2_2162 (N8436, N7114, N4661);
  and AND2_2167 (N8441, N7125, N4667);
  and AND2_2168 (N8442, N7136, N7125);
  and AND2_2171 (N8447, N7142, N4675);
  and AND2_2175 (N8451, N7149, N4678);
  and AND2_2178 (N8454, N4682, N7159);
  and AND2_2180 (N8456, N7170, N4687);
  and AND2_2222 (N8518, N7180, N7170);
  and AND2_2234 (N8545, N7346, N4757);
  and AND2_2238 (N8551, N7358, N4762);
  and AND2_2349 (N8818, N7609, N3122);
  and AND2_2359 (N8874, N6833, N7655);
  and AND2_2381 (N8960, N3375, N7852);
  and AND2_2477 (N9288, N367, N8326);
  and AND2_2490 (N9318, N8326, N6957);
  and AND2_2498 (N9332, N8405, N8412);
  and AND2_2500 (N9344, N8430, N8444);
  and AND2_2524 (N9385, N8430, N8497);
  and AND2_2537 (N9408, N8541, N8548);
  and AND2_2589 (N9526, N8943, N8421);
  and AND2_2594 (N9543, N8857, N8254);
  and AND2_2595 (N9551, N8871, N8288);
  and AND2_2599 (N9560, N8902, N8333);
  and AND2_2615 (N9585, N8405, N8956);
  and AND2_2616 (N9591, N8966, N8430);
  and AND2_2639 (N9618, N8541, N9035);
  and AND2_2689 (N9732, N9265, N8269);
  and AND2_2693 (N9736, N9265, N8262);
  and AND2_2700 (N9754, N8333, N9280);
  and AND2_2707 (N9767, N9280, N367);
  and AND2_2712 (N9775, N8333, N9307);
  and AND2_2735 (N9817, N9617, N9407);
  and AND2_2780 (N9932, N9575, N9773);
  and AND2_2781 (N9935, N9575, N9769);
  and AND2_2788 (N9949, N9608, N9375);
  and AND2_2849 (N10039, N9791, N8298);
  and AND2_2852 (N10042, N9758, N9385);
  and AND2_2856 (N10054, N9817, N9029);
  and AND2_2857 (N10055, N9786, N8394);
  and AND2_2859 (N10057, N9791, N8307);
  and AND2_2862 (N10060, N9758, N9344);
  and AND2_2881 (N10105, N9925, N9894);
  and AND2_2882 (N10106, N9925, N9895);
  and AND2_2883 (N10107, N9925, N9896);
  and AND2_2884 (N10108, N9925, N8253);
  and AND2_2895 (N10130, N9768, N9925);
  and AND2_2898 (N10133, N9932, N8898);
  and AND2_2904 (N10139, N9785, N10053);
  and AND2_2940 (N10230, N9768, N10131);
  and AND2_2956 (N10266, N10026, N10124);
  and AND2_2957 (N10267, N10028, N10124);
  and AND2_2958 (N10268, N9742, N10124);
  and AND2_2959 (N10269, N6923, N10124);
  and AND2_2967 (N10281, N10141, N5683);
  and AND2_2968 (N10282, N6784, N10141);
  and AND2_2973 (N10290, N10148, N5856);
  and AND2_2974 (N10291, N6881, N10148);
  and AND2_2975 (N10292, N8898, N10124);
  and AND2_2979 (N10296, N8959, N10234);
  and AND2_3014 (N10354, N8857, N10270);
  and AND2_3021 (N10391, N9582, N10295);
  and AND2_3042 (N10451, N10296, N4193);
  and AND2_3068 (N10546, N5631, N10450);
  and AND2_3070 (N10548, N10391, N8950);
  and AND2_3071 (N10549, N5165, N10367);
  and AND2_3073 (N10551, N10354, N3126);
  and AND2_3075 (N10553, N10375, N9539);
  and AND2_3076 (N10554, N10375, N9540);
  and AND2_3077 (N10555, N10375, N9541);
  and AND2_3078 (N10556, N10375, N6761);
  and AND2_3103 (N10587, N10367, N5735);
  and AND2_3104 (N10588, N10367, N3135);
  and AND2_3109 (N10597, N10381, N7180);
  and AND2_3110 (N10598, N8444, N10381);
  and AND2_3118 (N10629, N9733, N10547);
  and AND2_3119 (N10631, N5165, N10550);
  and AND2_3162 (N10705, N3126, N10583);
  and AND2_3164 (N10707, N9737, N10589);
  and AND2_3165 (N10708, N9738, N10589);
  and AND2_3166 (N10709, N9243, N10589);
  and AND2_3167 (N10710, N5850, N10589);
  and AND2_3179 (N10730, N5178, N10583);
  and AND2_3180 (N10731, N2523, N10583);
  and AND2_3197 (N10765, N10652, N9890);
  and AND2_3198 (N10766, N10652, N9891);
  and AND2_3199 (N10767, N10652, N9892);
  and AND2_3200 (N10768, N10652, N8252);
  and AND2_3246 (N10864, N10023, N10784);
  and AND2_3247 (N10865, N10024, N10784);
  and AND2_3248 (N10866, N9739, N10784);
  and AND2_3249 (N10867, N7136, N10784);
  and AND2_3466 (N11278, N10116, N11260);
  and AND2_3468 (N11280, N10119, N11262);
  and AND2_3474 (N11288, N11277, N10479);
  and AND2_3475 (N11289, N11279, N10283);
  and AND2_3484 (N11298, N10301, N11293);
  and AND2_3488 (N11308, N11296, N1115);
  and AND2_3489 (N11309, N11297, N10497);
  and AND2_3494 (N11316, N367, N11307);
  and AND3_1752 (N6767, N5640, N5632, N3101);
  and AND3_1756 (N6771, N5654, N3107, N5640);
  and AND3_1763 (N6778, N5670, N5654, N3114);
  and AND3_1764 (N6779, N5683, N5654, N5670);
  and AND3_1794 (N6837, N5778, N5771, N3173);
  and AND3_1797 (N6840, N5789, N3178, N5778);
  and AND3_1798 (N6841, N5850, N5789, N5778);
  and AND3_1804 (N6849, N5807, N5799, N3189);
  and AND3_1808 (N6853, N5821, N3195, N5807);
  and AND3_1815 (N6860, N5837, N5821, N3202);
  and AND3_1816 (N6861, N5856, N5821, N5837);
  and AND3_2075 (N8280, N5740, N5736, N5744);
  and AND3_2076 (N8281, N6800, N6797, N5744);
  and AND3_2077 (N8282, N5751, N5747, N5755);
  and AND3_2078 (N8283, N6806, N6803, N5755);
  and AND3_2079 (N8284, N5762, N5758, N5766);
  and AND3_2080 (N8285, N6812, N6809, N5766);
  and AND3_2099 (N8338, N6901, N6894, N4549);
  and AND3_2102 (N8341, N6912, N4555, N6901);
  and AND3_2103 (N8342, N6923, N6912, N6901);
  and AND3_2110 (N8349, N6936, N6929, N4566);
  and AND3_2114 (N8353, N6946, N4570, N6936);
  and AND3_2117 (N8356, N6957, N6946, N5960);
  and AND3_2160 (N8434, N7114, N7107, N4661);
  and AND3_2163 (N8437, N7125, N4667, N7114);
  and AND3_2164 (N8438, N7136, N7125, N7114);
  and AND3_2172 (N8448, N7149, N7142, N4678);
  and AND3_2176 (N8452, N7159, N4682, N7149);
  and AND3_2179 (N8455, N7170, N7159, N4687);
  and AND3_2191 (N8483, N6083, N6079, N6087);
  and AND3_2192 (N8484, N7191, N7188, N6087);
  and AND3_2217 (N8513, N7180, N7159, N7170);
  and AND3_2231 (N8539, N6141, N6137, N6145);
  and AND3_2232 (N8540, N7337, N7334, N6145);
  and AND3_2251 (N8578, N6170, N6166, N6174);
  and AND3_2252 (N8579, N7381, N7378, N6174);
  and AND3_2352 (N8861, N6797, N5740, N8274);
  and AND3_2353 (N8862, N5736, N6800, N8274);
  and AND3_2354 (N8863, N6803, N5751, N8276);
  and AND3_2355 (N8864, N5747, N6806, N8276);
  and AND3_2356 (N8865, N6809, N5762, N8278);
  and AND3_2357 (N8866, N5758, N6812, N8278);
  and AND3_2384 (N8991, N7188, N6083, N8469);
  and AND3_2385 (N8992, N6079, N7191, N8469);
  and AND3_2390 (N9024, N7334, N6141, N8537);
  and AND3_2391 (N9025, N6137, N7337, N8537);
  and AND3_2394 (N9053, N7378, N6170, N8564);
  and AND3_2395 (N9054, N6166, N7381, N8564);
  and AND3_2476 (N9287, N367, N8326, N6957);
  and AND3_2489 (N9315, N8326, N6946, N6957);
  and AND3_2515 (N9369, N7198, N7194, N7202);
  and AND3_2516 (N9370, N8460, N8457, N7202);
  and AND3_2517 (N9371, N7209, N7205, N7213);
  and AND3_2518 (N9372, N8466, N8463, N7213);
  and AND3_2529 (N9396, N7318, N7314, N7322);
  and AND3_2530 (N9397, N8522, N8519, N7322);
  and AND3_2531 (N9398, N6131, N6127, N7331);
  and AND3_2532 (N9399, N7328, N7325, N7331);
  and AND3_2545 (N9419, N7387, N6177, N7391);
  and AND3_2546 (N9420, N8555, N7384, N7391);
  and AND3_2547 (N9421, N7398, N7394, N7402);
  and AND3_2548 (N9422, N8561, N8558, N7402);
  and AND3_2627 (N9602, N8457, N7198, N9363);
  and AND3_2628 (N9603, N7194, N8460, N9363);
  and AND3_2629 (N9604, N8463, N7209, N9365);
  and AND3_2630 (N9605, N7205, N8466, N9365);
  and AND3_2633 (N9612, N8519, N7318, N9392);
  and AND3_2634 (N9613, N7314, N8522, N9392);
  and AND3_2635 (N9614, N7325, N6131, N9394);
  and AND3_2636 (N9615, N6127, N7328, N9394);
  and AND3_2640 (N9621, N7384, N7387, N9413);
  and AND3_2641 (N9622, N6177, N8555, N9413);
  and AND3_2642 (N9623, N8558, N7398, N9415);
  and AND3_2643 (N9624, N7394, N8561, N9415);
  and AND3_2827 (N10013, N9791, N8307, N8269);
  and AND3_2830 (N10016, N9786, N8394, N8421);
  and AND3_2834 (N10020, N9791, N8298, N8262);
  and AND3_2850 (N10040, N9758, N9385, N8298);
  and AND3_2853 (N10043, N367, N9775, N9385);
  and AND3_2858 (N10056, N9820, N9332, N8394);
  and AND3_2860 (N10058, N9758, N9344, N8307);
  and AND3_2863 (N10061, N367, N9754, N9344);
  and AND3_2966 (N10280, N10141, N5683, N5670);
  and AND3_2972 (N10289, N10148, N5856, N5837);
  and AND3_3099 (N10577, N10399, N10402, N10388);
  and AND3_3100 (N10581, N10360, N9543, N10116);
  and AND3_3101 (N10582, N10357, N9905, N10116);
  and AND3_3108 (N10596, N10381, N7180, N7170);
  and AND3_3130 (N10647, N886, N887, N10577);
  and AND3_3131 (N10648, N10360, N8857, N10479);
  and AND3_3132 (N10649, N10357, N7609, N10479);
  and AND3_3402 (N11152, N11103, N8871, N10283);
  and AND3_3403 (N11153, N11100, N7655, N10283);
  and AND3_3404 (N11154, N11103, N9551, N10119);
  and AND3_3405 (N11155, N11100, N9917, N10119);
  and AND3_3433 (N11222, N11159, N9575, N1115);
  and AND3_3434 (N11223, N11156, N8902, N1115);
  and AND3_3435 (N11224, N11159, N9935, N367);
  and AND3_3436 (N11225, N11156, N10132, N367);
  and AND3_3437 (N11226, N11165, N9608, N10497);
  and AND3_3438 (N11227, N11162, N8966, N10497);
  and AND3_3439 (N11228, N11165, N9949, N10301);
  and AND3_3440 (N11229, N11162, N10160, N10301);
  and AND4_11 (N494, N162, N172, N188, N199);
  and AND4_21 (N528, N150, N184, N228, N240);
  and AND4_41 (N575, N183, N182, N185, N186);
  and AND4_42 (N578, N210, N152, N218, N230);
  and AND4_1753 (N6768, N5654, N5632, N3107, N5640);
  and AND4_1757 (N6772, N5670, N5654, N3114, N5640);
  and AND4_1758 (N6773, N5683, N5654, N5640, N5670);
  and AND4_1792 (N6833, N5850, N5789, N5778, N5771);
  and AND4_1795 (N6838, N5789, N5771, N3178, N5778);
  and AND4_1805 (N6850, N5821, N5799, N3195, N5807);
  and AND4_1809 (N6854, N5837, N5821, N3202, N5807);
  and AND4_1810 (N6855, N5856, N5821, N5807, N5837);
  and AND4_1866 (N7057, N6021, N6000, N5996, N5991);
  and AND4_1869 (N7062, N6000, N5991, N3364, N5996);
  and AND4_1873 (N7066, N6014, N6003, N3368, N6009);
  and AND4_1887 (N7105, N6052, N6041, N3373, N6047);
  and AND4_2097 (N8333, N6901, N6923, N6912, N6894);
  and AND4_2100 (N8339, N6912, N6894, N4555, N6901);
  and AND4_2111 (N8350, N6946, N6929, N4570, N6936);
  and AND4_2115 (N8354, N6957, N6946, N5960, N6936);
  and AND4_2148 (N8405, N7098, N7077, N7073, N7068);
  and AND4_2151 (N8411, N7077, N7068, N4635, N7073);
  and AND4_2155 (N8417, N7091, N7080, N4640, N7086);
  and AND4_2158 (N8430, N7114, N7136, N7125, N7107);
  and AND4_2161 (N8435, N7125, N7107, N4667, N7114);
  and AND4_2173 (N8449, N7159, N7142, N4682, N7149);
  and AND4_2177 (N8453, N7170, N7159, N4687, N7149);
  and AND4_2211 (N8507, N7180, N7159, N7149, N7170);
  and AND4_2233 (N8541, N7376, N7355, N7351, N7346);
  and AND4_2236 (N8547, N7355, N7346, N4759, N7351);
  and AND4_2240 (N8553, N7369, N7358, N4766, N7364);
  and AND4_2475 (N9286, N367, N8326, N6946, N6957);
  and AND4_2488 (N9314, N8326, N6946, N6936, N6957);
  and AND4_2717 (N9790, N89, N9408, N9332, N8394);
  and AND4_2828 (N10014, N9758, N9344, N8307, N8269);
  and AND4_2831 (N10017, N9820, N9332, N8394, N8421);
  and AND4_2835 (N10021, N9758, N9385, N8298, N8262);
  and AND4_2851 (N10041, N367, N9775, N9385, N8298);
  and AND4_2861 (N10059, N367, N9754, N9344, N8307);
  and AND4_2965 (N10279, N10141, N5683, N5654, N5670);
  and AND4_2971 (N10288, N10148, N5856, N5821, N5837);
  and AND4_3020 (N10388, N10114, N10134, N10293, N10294);
  and AND4_3022 (N10399, N10113, N10115, N10299, N10300);
  and AND4_3023 (N10402, N10155, N10161, N10306, N10307);
  and AND4_3107 (N10595, N10381, N7180, N7159, N7170);
  nand NAND2_53 (N628, N12, N9);
  nand NAND2_72 (N700, N382, N267);
  nand NAND2_108 (N881, N467, N585);
  nand NAND2_119 (N1029, N382, N705);
  nand NAND2_121 (N1110, N242, N585);
  nand NAND2_393 (N2107, N38, N1821);
  nand NAND2_394 (N2108, N700, N1822);
  nand NAND2_396 (N2111, N957, N1822);
  nand NAND2_403 (N2172, N1029, N1822);
  nand NAND2_425 (N2257, N2107, N2108);
  nand NAND2_427 (N2268, N38, N688);
  nand NAND2_484 (N2355, N38, N2171);
  nand NAND2_486 (N2357, N1222, N1822);
  nand NAND2_558 (N2523, N2268, N2111);
  nand NAND2_578 (N2650, N2355, N2172);
  nand NAND2_579 (N2653, N38, N1028);
  nand NAND2_644 (N2988, N2653, N2357);
  nand NAND2_915 (N3953, N2257, N2117);
  nand NAND2_917 (N3955, N2257, N2537);
  nand NAND2_925 (N4326, N2769, N3551);
  nand NAND2_926 (N4327, N2766, N3552);
  nand NAND2_927 (N4333, N2775, N3569);
  nand NAND2_928 (N4334, N2772, N3570);
  nand NAND2_929 (N4411, N2787, N3781);
  nand NAND2_930 (N4412, N2784, N3782);
  nand NAND2_931 (N4463, N2644, N260);
  nand NAND2_933 (N4465, N2638, N257);
  nand NAND2_935 (N4467, N2632, N106);
  nand NAND2_937 (N4469, N2626, N254);
  nand NAND2_939 (N4471, N2619, N251);
  nand NAND2_955 (N4487, N1708, N3954);
  nand NAND2_956 (N4488, N1537, N3954);
  nand NAND2_958 (N4490, N2619, N628);
  nand NAND2_964 (N4496, N628, N2441);
  nand NAND2_970 (N4502, N2554, N3167);
  nand NAND2_975 (N4507, N2508, N303);
  nand NAND2_977 (N4509, N2502, N299);
  nand NAND2_979 (N4511, N2496, N296);
  nand NAND2_981 (N4513, N2482, N289);
  nand NAND2_983 (N4515, N2573, N286);
  nand NAND2_985 (N4517, N2567, N283);
  nand NAND2_987 (N4519, N2561, N280);
  nand NAND2_989 (N4521, N2488, N293);
  nand NAND2_991 (N4523, N2554, N277);
  nand NAND2_1083 (N4694, N2654, N3380);
  nand NAND2_1102 (N4746, N2604, N3452);
  nand NAND2_1107 (N4751, N2538, N3453);
  nand NAND2_1127 (N4776, N2729, N3486);
  nand NAND2_1146 (N4803, N4326, N4327);
  nand NAND2_1147 (N4806, N4333, N4334);
  nand NAND2_1212 (N4997, N4411, N4412);
  nand NAND2_1276 (N5165, N3507, N4473);
  nand NAND2_1278 (N5167, N666, N4464);
  nand NAND2_1279 (N5168, N660, N4466);
  nand NAND2_1280 (N5169, N674, N4468);
  nand NAND2_1281 (N5170, N651, N4470);
  nand NAND2_1282 (N5171, N644, N4472);
  nand NAND2_1288 (N5177, N3953, N4487);
  nand NAND2_1289 (N5178, N3955, N4488);
  nand NAND2_1290 (N5179, N3073, N4472);
  nand NAND2_1291 (N5180, N2626, N4468);
  nand NAND2_1292 (N5181, N2632, N4470);
  nand NAND2_1293 (N5182, N2638, N4464);
  nand NAND2_1294 (N5183, N2644, N4466);
  nand NAND2_1295 (N5184, N3080, N3073);
  nand NAND2_1296 (N5185, N2446, N4497);
  nand NAND2_1297 (N5186, N2450, N4498);
  nand NAND2_1298 (N5187, N2454, N4499);
  nand NAND2_1299 (N5188, N2458, N4500);
  nand NAND2_1300 (N5189, N2778, N4501);
  nand NAND2_1301 (N5190, N2561, N4503);
  nand NAND2_1302 (N5191, N2567, N4504);
  nand NAND2_1303 (N5192, N2573, N4505);
  nand NAND2_1304 (N5193, N2482, N4506);
  nand NAND2_1305 (N5196, N609, N4508);
  nand NAND2_1306 (N5197, N604, N4510);
  nand NAND2_1307 (N5198, N742, N4512);
  nand NAND2_1308 (N5199, N599, N4505);
  nand NAND2_1309 (N5200, N727, N4506);
  nand NAND2_1310 (N5201, N721, N4503);
  nand NAND2_1311 (N5202, N715, N4504);
  nand NAND2_1312 (N5203, N734, N4522);
  nand NAND2_1313 (N5204, N708, N4501);
  nand NAND2_1323 (N5283, N2478, N4611);
  nand NAND2_1324 (N5284, N2761, N4612);
  nand NAND2_1325 (N5285, N2474, N4613);
  nand NAND2_1326 (N5286, N2757, N4614);
  nand NAND2_1327 (N5287, N2470, N4615);
  nand NAND2_1328 (N5288, N2753, N4616);
  nand NAND2_1329 (N5289, N2462, N4617);
  nand NAND2_1330 (N5290, N2745, N4618);
  nand NAND2_1331 (N5291, N2550, N4619);
  nand NAND2_1332 (N5292, N2741, N4620);
  nand NAND2_1333 (N5293, N2546, N4621);
  nand NAND2_1334 (N5294, N2737, N4622);
  nand NAND2_1335 (N5295, N2542, N4623);
  nand NAND2_1336 (N5296, N2733, N4624);
  nand NAND2_1337 (N5297, N2466, N4625);
  nand NAND2_1338 (N5298, N2749, N4626);
  nand NAND2_1339 (N5299, N2538, N4627);
  nand NAND2_1340 (N5300, N2729, N4628);
  nand NAND2_1341 (N5314, N2458, N4643);
  nand NAND2_1342 (N5315, N2670, N4499);
  nand NAND2_1343 (N5316, N2454, N4645);
  nand NAND2_1344 (N5317, N2666, N4500);
  nand NAND2_1345 (N5318, N2450, N4647);
  nand NAND2_1346 (N5319, N2662, N4497);
  nand NAND2_1347 (N5320, N2446, N4649);
  nand NAND2_1348 (N5321, N2658, N4498);
  nand NAND2_1349 (N5322, N628, N4651);
  nand NAND2_1350 (N5323, N2654, N3073);
  nand NAND2_1352 (N5363, N2781, N4651);
  nand NAND2_1353 (N5364, N2658, N4647);
  nand NAND2_1354 (N5365, N2662, N4649);
  nand NAND2_1355 (N5366, N2666, N4643);
  nand NAND2_1356 (N5367, N2670, N4645);
  nand NAND2_1357 (N5425, N2790, N4745);
  nand NAND2_1358 (N5426, N2607, N4747);
  nand NAND2_1359 (N5427, N2611, N4748);
  nand NAND2_1360 (N5429, N2793, N4628);
  nand NAND2_1361 (N5430, N2542, N4622);
  nand NAND2_1362 (N5431, N2546, N4624);
  nand NAND2_1363 (N5432, N2550, N4618);
  nand NAND2_1364 (N5433, N2462, N4620);
  nand NAND2_1365 (N5451, N2796, N4627);
  nand NAND2_1366 (N5452, N2733, N4621);
  nand NAND2_1367 (N5453, N2737, N4623);
  nand NAND2_1368 (N5454, N2741, N4617);
  nand NAND2_1369 (N5455, N2745, N4619);
  nand NAND2_1370 (N5456, N3888, N4781);
  nand NAND2_1371 (N5457, N3885, N4782);
  nand NAND2_1373 (N5474, N2488, N4512);
  nand NAND2_1374 (N5475, N2496, N4522);
  nand NAND2_1375 (N5476, N2502, N4508);
  nand NAND2_1376 (N5477, N2508, N4510);
  nand NAND2_1377 (N5571, N2692, N4633);
  nand NAND2_1378 (N5572, N2696, N4642);
  nand NAND2_1379 (N5573, N2700, N4629);
  nand NAND2_1380 (N5574, N2704, N4631);
  nand NAND2_1381 (N5584, N2466, N4616);
  nand NAND2_1382 (N5585, N2470, N4626);
  nand NAND2_1383 (N5586, N2474, N4612);
  nand NAND2_1384 (N5587, N2478, N4614);
  nand NAND2_1385 (N5602, N2749, N4615);
  nand NAND2_1386 (N5603, N2753, N4625);
  nand NAND2_1387 (N5604, N2757, N4611);
  nand NAND2_1388 (N5605, N2761, N4613);
  nand NAND2_1389 (N5631, N5324, N4653);
  nand NAND2_1390 (N5632, N4463, N5167);
  nand NAND2_1391 (N5640, N4465, N5168);
  nand NAND2_1392 (N5654, N4467, N5169);
  nand NAND2_1393 (N5670, N4469, N5170);
  nand NAND2_1394 (N5683, N4471, N5171);
  nand NAND2_1401 (N5736, N5179, N4490);
  nand NAND2_1402 (N5740, N5180, N5181);
  nand NAND2_1403 (N5744, N5182, N5183);
  nand NAND2_1404 (N5747, N5184, N4496);
  nand NAND2_1405 (N5751, N5185, N5186);
  nand NAND2_1406 (N5755, N5187, N5188);
  nand NAND2_1407 (N5758, N5189, N4502);
  nand NAND2_1408 (N5762, N5190, N5191);
  nand NAND2_1409 (N5766, N5192, N5193);
  nand NAND2_1412 (N5771, N4507, N5196);
  nand NAND2_1413 (N5778, N4509, N5197);
  nand NAND2_1414 (N5789, N4511, N5198);
  nand NAND2_1415 (N5799, N4513, N5199);
  nand NAND2_1416 (N5807, N4515, N5200);
  nand NAND2_1417 (N5821, N4517, N5201);
  nand NAND2_1418 (N5837, N4519, N5202);
  nand NAND2_1419 (N5850, N4521, N5203);
  nand NAND2_1420 (N5856, N4523, N5204);
  nand NAND2_1431 (N5944, N3293, N334);
  nand NAND2_1433 (N5946, N3287, N331);
  nand NAND2_1435 (N5948, N3281, N328);
  nand NAND2_1437 (N5950, N3273, N325);
  nand NAND2_1439 (N5952, N3267, N322);
  nand NAND2_1441 (N5954, N3355, N319);
  nand NAND2_1443 (N5956, N3349, N316);
  nand NAND2_1445 (N5958, N3343, N313);
  nand NAND2_1466 (N5991, N5283, N5284);
  nand NAND2_1467 (N5996, N5285, N5286);
  nand NAND2_1468 (N6000, N5287, N5288);
  nand NAND2_1469 (N6003, N5289, N5290);
  nand NAND2_1470 (N6009, N5291, N5292);
  nand NAND2_1471 (N6014, N5293, N5294);
  nand NAND2_1472 (N6018, N5295, N5296);
  nand NAND2_1473 (N6021, N5297, N5298);
  nand NAND2_1474 (N6022, N5299, N5300);
  nand NAND2_1476 (N6024, N3448, N4629);
  nand NAND2_1478 (N6026, N3444, N4631);
  nand NAND2_1480 (N6028, N3440, N4633);
  nand NAND2_1482 (N6030, N3432, N4636);
  nand NAND2_1490 (N6038, N3436, N4642);
  nand NAND2_1493 (N6041, N5314, N5315);
  nand NAND2_1494 (N6047, N5316, N5317);
  nand NAND2_1495 (N6052, N5318, N5319);
  nand NAND2_1496 (N6056, N5320, N5321);
  nand NAND2_1497 (N6059, N5322, N5323);
  nand NAND2_1498 (N6060, N3410, N364);
  nand NAND2_1500 (N6062, N3404, N361);
  nand NAND2_1502 (N6064, N3398, N358);
  nand NAND2_1504 (N6066, N3390, N355);
  nand NAND2_1506 (N6068, N3384, N352);
  nand NAND2_1508 (N6070, N3334, N349);
  nand NAND2_1510 (N6072, N3328, N346);
  nand NAND2_1512 (N6074, N3322, N343);
  nand NAND2_1514 (N6076, N3315, N340);
  nand NAND2_1517 (N6079, N5363, N4694);
  nand NAND2_1518 (N6083, N5364, N5365);
  nand NAND2_1519 (N6087, N5366, N5367);
  nand NAND2_1521 (N6091, N3315, N4699);
  nand NAND2_1527 (N6097, N3340, N4700);
  nand NAND2_1552 (N6122, N3299, N4743);
  nand NAND2_1555 (N6125, N3311, N4636);
  nand NAND2_1557 (N6127, N5425, N4746);
  nand NAND2_1558 (N6131, N5426, N5427);
  nand NAND2_1560 (N6136, N3247, N4749);
  nand NAND2_1561 (N6137, N5429, N4751);
  nand NAND2_1562 (N6141, N5430, N5431);
  nand NAND2_1563 (N6145, N5432, N5433);
  nand NAND2_1573 (N6157, N3462, N4749);
  nand NAND2_1575 (N6159, N3458, N4747);
  nand NAND2_1577 (N6161, N3454, N4748);
  nand NAND2_1580 (N6164, N3381, N4768);
  nand NAND2_1582 (N6166, N5451, N4776);
  nand NAND2_1583 (N6170, N5452, N5453);
  nand NAND2_1584 (N6174, N5454, N5455);
  nand NAND2_1585 (N6177, N5456, N5457);
  nand NAND2_1591 (N6186, N3416, N4783);
  nand NAND2_1597 (N6192, N4784, N2117);
  nand NAND2_1599 (N6194, N3507, N2537);
  nand NAND2_1601 (N6196, N5476, N5477);
  nand NAND2_1602 (N6199, N5474, N5475);
  nand NAND2_1628 (N6243, N5573, N5574);
  nand NAND2_1629 (N6246, N5571, N5572);
  nand NAND2_1630 (N6249, N5586, N5587);
  nand NAND2_1631 (N6252, N5584, N5585);
  nand NAND2_1640 (N6263, N5604, N5605);
  nand NAND2_1641 (N6266, N5602, N5603);
  nand NAND2_1642 (N6540, N806, N5945);
  nand NAND2_1643 (N6541, N800, N5947);
  nand NAND2_1644 (N6542, N794, N5949);
  nand NAND2_1645 (N6543, N786, N5951);
  nand NAND2_1646 (N6544, N780, N5953);
  nand NAND2_1647 (N6545, N774, N5955);
  nand NAND2_1648 (N6546, N768, N5957);
  nand NAND2_1649 (N6547, N762, N5959);
  nand NAND2_1658 (N6594, N2704, N6023);
  nand NAND2_1659 (N6595, N2700, N6025);
  nand NAND2_1660 (N6596, N2696, N6027);
  nand NAND2_1661 (N6597, N2688, N6029);
  nand NAND2_1662 (N6598, N3311, N6031);
  nand NAND2_1663 (N6599, N3428, N6032);
  nand NAND2_1664 (N6600, N3307, N6033);
  nand NAND2_1665 (N6601, N3424, N6034);
  nand NAND2_1666 (N6602, N3303, N6035);
  nand NAND2_1667 (N6603, N3420, N6036);
  nand NAND2_1668 (N6604, N2692, N6037);
  nand NAND2_1669 (N6605, N3299, N6039);
  nand NAND2_1670 (N6606, N3416, N6040);
  nand NAND2_1671 (N6621, N865, N6061);
  nand NAND2_1672 (N6622, N859, N6063);
  nand NAND2_1673 (N6623, N853, N6065);
  nand NAND2_1674 (N6624, N845, N6067);
  nand NAND2_1675 (N6625, N839, N6069);
  nand NAND2_1676 (N6626, N833, N6071);
  nand NAND2_1677 (N6627, N827, N6073);
  nand NAND2_1678 (N6628, N821, N6075);
  nand NAND2_1679 (N6629, N814, N6077);
  nand NAND2_1680 (N6639, N3783, N6077);
  nand NAND2_1681 (N6640, N3322, N6073);
  nand NAND2_1682 (N6641, N3328, N6075);
  nand NAND2_1683 (N6642, N3334, N6069);
  nand NAND2_1684 (N6643, N3384, N6071);
  nand NAND2_1685 (N6644, N3786, N6096);
  nand NAND2_1686 (N6645, N3343, N5957);
  nand NAND2_1687 (N6646, N3349, N5959);
  nand NAND2_1688 (N6647, N3355, N5953);
  nand NAND2_1689 (N6648, N3267, N5955);
  nand NAND2_1699 (N6658, N3789, N6040);
  nand NAND2_1700 (N6659, N3303, N6034);
  nand NAND2_1701 (N6660, N3307, N6036);
  nand NAND2_1702 (N6661, N2688, N6032);
  nand NAND2_1703 (N6668, N2615, N6135);
  nand NAND2_1704 (N6677, N3263, N6148);
  nand NAND2_1705 (N6678, N3482, N6149);
  nand NAND2_1706 (N6679, N3259, N6150);
  nand NAND2_1707 (N6680, N3478, N6151);
  nand NAND2_1708 (N6681, N3255, N6152);
  nand NAND2_1709 (N6682, N3474, N6153);
  nand NAND2_1710 (N6683, N3247, N6154);
  nand NAND2_1711 (N6684, N3466, N6135);
  nand NAND2_1712 (N6685, N2615, N6156);
  nand NAND2_1713 (N6686, N2611, N6158);
  nand NAND2_1714 (N6687, N2607, N6160);
  nand NAND2_1715 (N6688, N3251, N6162);
  nand NAND2_1716 (N6689, N3470, N6163);
  nand NAND2_1717 (N6690, N2680, N6165);
  nand NAND2_1718 (N6702, N3454, N6158);
  nand NAND2_1719 (N6703, N3458, N6160);
  nand NAND2_1720 (N6704, N3462, N6154);
  nand NAND2_1721 (N6705, N3466, N6156);
  nand NAND2_1722 (N6706, N3891, N6039);
  nand NAND2_1723 (N6707, N3420, N6033);
  nand NAND2_1724 (N6708, N3424, N6035);
  nand NAND2_1725 (N6709, N3428, N6029);
  nand NAND2_1726 (N6710, N3432, N6031);
  nand NAND2_1727 (N6711, N1708, N6191);
  nand NAND2_1728 (N6712, N1537, N3126);
  nand NAND2_1729 (N6729, N3390, N6065);
  nand NAND2_1730 (N6730, N3398, N6067);
  nand NAND2_1731 (N6731, N3404, N6061);
  nand NAND2_1732 (N6732, N3410, N6063);
  nand NAND2_1733 (N6733, N3273, N5949);
  nand NAND2_1734 (N6734, N3281, N5951);
  nand NAND2_1735 (N6735, N3287, N5945);
  nand NAND2_1736 (N6736, N3293, N5947);
  nand NAND2_1737 (N6741, N3251, N6153);
  nand NAND2_1738 (N6742, N3255, N6163);
  nand NAND2_1739 (N6743, N3259, N6149);
  nand NAND2_1740 (N6744, N3263, N6151);
  nand NAND2_1741 (N6751, N3470, N6152);
  nand NAND2_1742 (N6752, N3474, N6162);
  nand NAND2_1743 (N6753, N3478, N6148);
  nand NAND2_1744 (N6754, N3482, N6150);
  nand NAND2_1745 (N6755, N3436, N6027);
  nand NAND2_1746 (N6756, N3440, N6037);
  nand NAND2_1747 (N6757, N3444, N6023);
  nand NAND2_1748 (N6758, N3448, N6025);
  nand NAND2_1845 (N6894, N5944, N6540);
  nand NAND2_1846 (N6901, N5946, N6541);
  nand NAND2_1847 (N6912, N5948, N6542);
  nand NAND2_1848 (N6923, N5950, N6543);
  nand NAND2_1849 (N6929, N5952, N6544);
  nand NAND2_1850 (N6936, N5954, N6545);
  nand NAND2_1851 (N6946, N5956, N6546);
  nand NAND2_1852 (N6957, N5958, N6547);
  nand NAND2_1853 (N6967, N4769, N4575);
  nand NAND2_1875 (N7068, N6594, N6024);
  nand NAND2_1876 (N7073, N6595, N6026);
  nand NAND2_1877 (N7077, N6596, N6028);
  nand NAND2_1878 (N7080, N6597, N6030);
  nand NAND2_1879 (N7086, N6598, N6599);
  nand NAND2_1880 (N7091, N6600, N6601);
  nand NAND2_1881 (N7095, N6602, N6603);
  nand NAND2_1882 (N7098, N6604, N6038);
  nand NAND2_1883 (N7099, N6605, N6606);
  nand NAND2_1889 (N7107, N6060, N6621);
  nand NAND2_1890 (N7114, N6062, N6622);
  nand NAND2_1891 (N7125, N6064, N6623);
  nand NAND2_1892 (N7136, N6066, N6624);
  nand NAND2_1893 (N7142, N6068, N6625);
  nand NAND2_1894 (N7149, N6070, N6626);
  nand NAND2_1895 (N7159, N6072, N6627);
  nand NAND2_1896 (N7170, N6074, N6628);
  nand NAND2_1897 (N7180, N6076, N6629);
  nand NAND2_1901 (N7194, N6639, N6091);
  nand NAND2_1902 (N7198, N6640, N6641);
  nand NAND2_1903 (N7202, N6642, N6643);
  nand NAND2_1904 (N7205, N6644, N6097);
  nand NAND2_1905 (N7209, N6645, N6646);
  nand NAND2_1906 (N7213, N6647, N6648);
  nand NAND2_1918 (N7314, N6658, N6122);
  nand NAND2_1919 (N7318, N6659, N6660);
  nand NAND2_1920 (N7322, N6125, N6661);
  nand NAND2_1923 (N7331, N6668, N6136);
  nand NAND2_1928 (N7346, N6677, N6678);
  nand NAND2_1929 (N7351, N6679, N6680);
  nand NAND2_1930 (N7355, N6681, N6682);
  nand NAND2_1931 (N7358, N6683, N6684);
  nand NAND2_1932 (N7364, N6685, N6157);
  nand NAND2_1933 (N7369, N6686, N6159);
  nand NAND2_1934 (N7373, N6687, N6161);
  nand NAND2_1935 (N7376, N6688, N6689);
  nand NAND2_1936 (N7377, N6164, N6690);
  nand NAND2_1940 (N7387, N6702, N6703);
  nand NAND2_1941 (N7391, N6704, N6705);
  nand NAND2_1942 (N7394, N6706, N6186);
  nand NAND2_1943 (N7398, N6707, N6708);
  nand NAND2_1944 (N7402, N6709, N6710);
  nand NAND2_1957 (N7441, N6192, N6711);
  nand NAND2_1958 (N7444, N6194, N6712);
  nand NAND2_2002 (N7560, N6731, N6732);
  nand NAND2_2003 (N7563, N6729, N6730);
  nand NAND2_2004 (N7566, N6735, N6736);
  nand NAND2_2005 (N7569, N6733, N6734);
  nand NAND2_2008 (N7574, N6743, N6744);
  nand NAND2_2009 (N7577, N6741, N6742);
  nand NAND2_2012 (N7582, N6753, N6754);
  nand NAND2_2013 (N7585, N6751, N6752);
  nand NAND2_2014 (N7588, N6757, N6758);
  nand NAND2_2015 (N7591, N6755, N6756);
  nand NAND2_2025 (N7744, N2674, N6968);
  nand NAND2_2034 (N8144, N6199, N7477);
  nand NAND2_2035 (N8145, N6196, N7478);
  nand NAND2_2046 (N8216, N6252, N7556);
  nand NAND2_2047 (N8217, N6249, N7557);
  nand NAND2_2048 (N8218, N6246, N7558);
  nand NAND2_2049 (N8219, N6243, N7559);
  nand NAND2_2050 (N8232, N6266, N7580);
  nand NAND2_2051 (N8233, N6263, N7581);
  nand NAND2_2092 (N8322, N5789, N4543);
  nand NAND2_2094 (N8324, N5789, N5943);
  nand NAND2_2096 (N8326, N6967, N7744);
  nand NAND2_2263 (N8608, N7441, N5469);
  nand NAND2_2265 (N8610, N7444, N3126);
  nand NAND2_2274 (N8627, N8144, N8145);
  nand NAND2_2312 (N8727, N8216, N8217);
  nand NAND2_2313 (N8730, N8218, N8219);
  nand NAND2_2344 (N8811, N8232, N8233);
  nand NAND2_2362 (N8880, N8146, N8315);
  nand NAND2_2364 (N8882, N8156, N8315);
  nand NAND2_2366 (N8884, N8204, N8294);
  nand NAND2_2368 (N8886, N8208, N8294);
  nand NAND2_2369 (N8887, N3625, N8323);
  nand NAND2_2370 (N8888, N3178, N8323);
  nand NAND2_2396 (N9064, N4303, N8607);
  nand NAND2_2397 (N9065, N3507, N8609);
  nand NAND2_2399 (N9067, N8114, N4795);
  nand NAND2_2403 (N9073, N8131, N6195);
  nand NAND2_2411 (N9088, N8166, N4813);
  nand NAND2_2415 (N9094, N8183, N6203);
  nand NAND2_2426 (N9159, N7577, N8733);
  nand NAND2_2427 (N9160, N7574, N8734);
  nand NAND2_2432 (N9179, N7563, N8753);
  nand NAND2_2433 (N9180, N7560, N8754);
  nand NAND2_2434 (N9181, N7569, N8755);
  nand NAND2_2435 (N9182, N7566, N8756);
  nand NAND2_2442 (N9234, N7591, N8814);
  nand NAND2_2443 (N9235, N7588, N8815);
  nand NAND2_2444 (N9236, N7585, N8816);
  nand NAND2_2445 (N9237, N7582, N8817);
  nand NAND2_2448 (N9243, N8324, N8888);
  nand NAND2_2467 (N9271, N5771, N8879);
  nand NAND2_2468 (N9272, N5771, N8881);
  nand NAND2_2469 (N9273, N5778, N8883);
  nand NAND2_2470 (N9274, N5778, N7650);
  nand NAND2_2471 (N9275, N8322, N8887);
  nand NAND2_2482 (N9297, N6912, N5966);
  nand NAND2_2484 (N9299, N6912, N6969);
  nand NAND2_2505 (N9359, N7125, N6078);
  nand NAND2_2507 (N9361, N7125, N7187);
  nand NAND2_2536 (N9407, N8548, N89);
  nand NAND2_2550 (N9426, N9064, N8608);
  nand NAND2_2551 (N9429, N9065, N8610);
  nand NAND2_2552 (N9432, N3515, N9066);
  nand NAND2_2553 (N9435, N3114, N9072);
  nand NAND2_2554 (N9442, N3628, N9087);
  nand NAND2_2555 (N9445, N3202, N9093);
  nand NAND2_2570 (N9478, N9159, N9160);
  nand NAND2_2571 (N9485, N9179, N9180);
  nand NAND2_2572 (N9488, N9181, N9182);
  nand NAND2_2587 (N9517, N9234, N9235);
  nand NAND2_2588 (N9520, N9236, N9237);
  nand NAND2_2591 (N9539, N9271, N8880);
  nand NAND2_2592 (N9540, N9273, N8884);
  nand NAND2_2596 (N9555, N9272, N8882);
  nand NAND2_2597 (N9556, N9274, N8886);
  nand NAND2_2601 (N9562, N9099, N9290);
  nand NAND2_2603 (N9564, N9103, N9290);
  nand NAND2_2605 (N9566, N9107, N9294);
  nand NAND2_2607 (N9568, N9111, N9294);
  nand NAND2_2608 (N9569, N4844, N9298);
  nand NAND2_2609 (N9570, N4555, N9298);
  nand NAND2_2618 (N9593, N9161, N9352);
  nand NAND2_2620 (N9595, N9165, N9352);
  nand NAND2_2622 (N9597, N9169, N9356);
  nand NAND2_2624 (N9599, N9173, N9356);
  nand NAND2_2625 (N9600, N4940, N9360);
  nand NAND2_2626 (N9601, N4667, N9360);
  nand NAND2_2648 (N9642, N9067, N9432);
  nand NAND2_2650 (N9646, N9073, N9435);
  nand NAND2_2652 (N9650, N9257, N9256);
  nand NAND2_2653 (N9653, N9259, N9258);
  nand NAND2_2654 (N9656, N9261, N9260);
  nand NAND2_2656 (N9660, N9079, N4543);
  nand NAND2_2658 (N9662, N8208, N5943);
  nand NAND2_2659 (N9663, N9088, N9442);
  nand NAND2_2661 (N9667, N9094, N9445);
  nand NAND2_2671 (N9691, N9146, N8717);
  nand NAND2_2674 (N9698, N9401, N9400);
  nand NAND2_2675 (N9702, N9368, N9367);
  nand NAND2_2681 (N9716, N9203, N6235);
  nand NAND2_2685 (N9722, N9220, N7573);
  nand NAND2_2688 (N9727, N9418, N9417);
  nand NAND2_2690 (N9733, N9581, N9326);
  nand NAND2_2696 (N9739, N9361, N9601);
  nand NAND2_2697 (N9740, N8326, N1115);
  nand NAND2_2699 (N9742, N9299, N9570);
  nand NAND2_2702 (N9762, N6894, N9561);
  nand NAND2_2703 (N9763, N6894, N9563);
  nand NAND2_2704 (N9764, N6901, N9565);
  nand NAND2_2705 (N9765, N6901, N8924);
  nand NAND2_2706 (N9766, N9297, N9569);
  nand NAND2_2708 (N9768, N9557, N9276);
  nand NAND2_2710 (N9773, N9307, N367);
  nand NAND2_2715 (N9785, N9616, N9402);
  nand NAND2_2719 (N9795, N7107, N9592);
  nand NAND2_2720 (N9796, N7107, N9594);
  nand NAND2_2721 (N9797, N7114, N9596);
  nand NAND2_2722 (N9798, N7114, N8996);
  nand NAND2_2723 (N9799, N9359, N9600);
  nand NAND2_2744 (N9836, N9426, N3135);
  nand NAND2_2746 (N9838, N9429, N3135);
  nand NAND2_2747 (N9846, N3625, N9659);
  nand NAND2_2748 (N9847, N3178, N7650);
  nand NAND2_2750 (N9863, N5960, N9690);
  nand NAND2_2752 (N9873, N5030, N9715);
  nand NAND2_2753 (N9876, N4687, N9721);
  nand NAND2_2754 (N9890, N9795, N9593);
  nand NAND2_2755 (N9891, N9797, N9597);
  nand NAND2_2757 (N9893, N367, N9741);
  nand NAND2_2758 (N9894, N9762, N9562);
  nand NAND2_2759 (N9895, N9764, N9566);
  nand NAND2_2762 (N9898, N9626, N9249);
  nand NAND2_2764 (N9900, N9629, N9250);
  nand NAND2_2766 (N9902, N9632, N9251);
  nand NAND2_2768 (N9904, N9635, N9252);
  nand NAND2_2771 (N9907, N9650, N5769);
  nand NAND2_2773 (N9909, N9653, N5770);
  nand NAND2_2775 (N9911, N9656, N9262);
  nand NAND2_2777 (N9923, N9763, N9564);
  nand NAND2_2778 (N9924, N9765, N9568);
  nand NAND2_2783 (N9939, N9698, N9323);
  nand NAND2_2784 (N9945, N9796, N9595);
  nand NAND2_2785 (N9946, N9798, N9599);
  nand NAND2_2787 (N9948, N9702, N6102);
  nand NAND2_2790 (N9954, N9727, N9412);
  nand NAND2_2791 (N9955, N2523, N9835);
  nand NAND2_2792 (N9956, N2523, N9837);
  nand NAND2_2794 (N9958, N9642, N9645);
  nand NAND2_2796 (N9960, N9646, N7613);
  nand NAND2_2797 (N9961, N9660, N9846);
  nand NAND2_2798 (N9964, N9662, N9847);
  nand NAND2_2800 (N9968, N9663, N9666);
  nand NAND2_2802 (N9970, N9667, N7659);
  nand NAND2_2804 (N9972, N9671, N5966);
  nand NAND2_2806 (N9974, N9111, N6969);
  nand NAND2_2808 (N9976, N9679, N7552);
  nand NAND2_2811 (N9979, N9691, N9863);
  nand NAND2_2813 (N9983, N9814, N9813);
  nand NAND2_2814 (N9986, N9816, N9815);
  nand NAND2_2815 (N9989, N9801, N9800);
  nand NAND2_2816 (N9992, N9803, N9802);
  nand NAND2_2818 (N9996, N9707, N6078);
  nand NAND2_2820 (N9998, N9173, N7187);
  nand NAND2_2821 (N9999, N9716, N9873);
  nand NAND2_2823 (N10003, N9722, N9876);
  nand NAND2_2825 (N10007, N9830, N9829);
  nand NAND2_2826 (N10010, N9828, N9827);
  nand NAND2_2839 (N10025, N9740, N9893);
  nand NAND2_2842 (N10032, N6929, N9897);
  nand NAND2_2843 (N10033, N6936, N9899);
  nand NAND2_2844 (N10034, N6946, N9901);
  nand NAND2_2845 (N10035, N6957, N9903);
  nand NAND2_2846 (N10036, N4803, N9906);
  nand NAND2_2847 (N10037, N4806, N9908);
  nand NAND2_2848 (N10038, N8627, N9910);
  nand NAND2_2854 (N10050, N8727, N9938);
  nand NAND2_2864 (N10062, N4997, N9947);
  nand NAND2_2865 (N10067, N8811, N9953);
  nand NAND2_2866 (N10070, N9955, N9836);
  nand NAND2_2867 (N10073, N9956, N9838);
  nand NAND2_2868 (N10076, N9068, N9957);
  nand NAND2_2869 (N10077, N9074, N9959);
  nand NAND2_2870 (N10082, N9089, N9967);
  nand NAND2_2871 (N10083, N9095, N9969);
  nand NAND2_2872 (N10084, N4844, N9971);
  nand NAND2_2873 (N10085, N4555, N8924);
  nand NAND2_2874 (N10086, N6217, N9975);
  nand NAND2_2875 (N10093, N4940, N9995);
  nand NAND2_2876 (N10094, N4667, N8996);
  nand NAND2_2885 (N10109, N10032, N9898);
  nand NAND2_2886 (N10110, N10033, N9900);
  nand NAND2_2887 (N10111, N10034, N9902);
  nand NAND2_2888 (N10112, N10035, N9904);
  nand NAND2_2889 (N10113, N10036, N9907);
  nand NAND2_2890 (N10114, N10037, N9909);
  nand NAND2_2891 (N10115, N10038, N9911);
  nand NAND2_2899 (N10134, N10050, N9939);
  nand NAND2_2901 (N10136, N9983, N9324);
  nand NAND2_2903 (N10138, N9986, N9784);
  nand NAND2_2908 (N10155, N10062, N9948);
  nand NAND2_2910 (N10157, N9989, N9805);
  nand NAND2_2912 (N10159, N9992, N9806);
  nand NAND2_2914 (N10161, N10067, N9954);
  nand NAND2_2916 (N10163, N10007, N9825);
  nand NAND2_2918 (N10165, N10010, N9826);
  nand NAND2_2919 (N10170, N10076, N9958);
  nand NAND2_2920 (N10173, N10077, N9960);
  nand NAND2_2922 (N10177, N9961, N8879);
  nand NAND2_2924 (N10179, N9964, N8881);
  nand NAND2_2925 (N10180, N10082, N9968);
  nand NAND2_2926 (N10183, N10083, N9970);
  nand NAND2_2927 (N10186, N9972, N10084);
  nand NAND2_2928 (N10189, N9974, N10085);
  nand NAND2_2929 (N10192, N9976, N10086);
  nand NAND2_2931 (N10196, N9979, N8931);
  nand NAND2_2932 (N10197, N9996, N10093);
  nand NAND2_2933 (N10200, N9998, N10094);
  nand NAND2_2935 (N10204, N9999, N10002);
  nand NAND2_2937 (N10206, N10003, N9005);
  nand NAND2_2938 (N10212, N10070, N3954);
  nand NAND2_2939 (N10213, N10073, N3954);
  nand NAND2_2941 (N10231, N8730, N10135);
  nand NAND2_2942 (N10232, N9478, N10137);
  nand NAND2_2944 (N10234, N7100, N10140);
  nand NAND2_2945 (N10237, N9485, N10156);
  nand NAND2_2946 (N10238, N9488, N10158);
  nand NAND2_2947 (N10239, N9517, N10162);
  nand NAND2_2948 (N10240, N9520, N10164);
  nand NAND2_2951 (N10247, N8146, N10176);
  nand NAND2_2952 (N10248, N8156, N10178);
  nand NAND2_2953 (N10259, N9692, N10195);
  nand NAND2_2954 (N10264, N9717, N10203);
  nand NAND2_2955 (N10265, N9723, N10205);
  nand NAND2_2960 (N10270, N6762, N10116);
  nand NAND2_2961 (N10271, N2257, N10241);
  nand NAND2_2962 (N10272, N2257, N10242);
  nand NAND2_2976 (N10293, N10231, N10136);
  nand NAND2_2977 (N10294, N10232, N10138);
  nand NAND2_2978 (N10295, N8412, N10233);
  nand NAND2_2980 (N10299, N10237, N10157);
  nand NAND2_2981 (N10300, N10238, N10159);
  nand NAND2_2983 (N10306, N10239, N10163);
  nand NAND2_2984 (N10307, N10240, N10165);
  nand NAND2_2988 (N10315, N10170, N9071);
  nand NAND2_2990 (N10317, N10173, N9077);
  nand NAND2_2991 (N10318, N10247, N10177);
  nand NAND2_2992 (N10321, N10248, N10179);
  nand NAND2_2994 (N10325, N10180, N9092);
  nand NAND2_2996 (N10327, N10183, N9098);
  nand NAND2_2998 (N10329, N10186, N9561);
  nand NAND2_3000 (N10331, N10189, N9563);
  nand NAND2_3002 (N10333, N10192, N9977);
  nand NAND2_3003 (N10334, N10259, N10196);
  nand NAND2_3005 (N10338, N10197, N9592);
  nand NAND2_3007 (N10340, N10200, N9594);
  nand NAND2_3008 (N10341, N10264, N10204);
  nand NAND2_3009 (N10344, N10265, N10206);
  nand NAND2_3015 (N10357, N10271, N10212);
  nand NAND2_3016 (N10360, N10272, N10213);
  nand NAND2_3032 (N10431, N8117, N10314);
  nand NAND2_3033 (N10432, N8134, N10316);
  nand NAND2_3034 (N10437, N8169, N10324);
  nand NAND2_3035 (N10438, N8186, N10326);
  nand NAND2_3036 (N10439, N9099, N10328);
  nand NAND2_3037 (N10440, N9103, N10330);
  nand NAND2_3038 (N10441, N9682, N10332);
  nand NAND2_3039 (N10444, N9161, N10337);
  nand NAND2_3040 (N10445, N9165, N10339);
  nand NAND2_3044 (N10456, N10148, N8242);
  nand NAND2_3046 (N10466, N10141, N8247);
  nand NAND2_3049 (N10509, N10431, N10315);
  nand NAND2_3050 (N10512, N10432, N10317);
  nand NAND2_3052 (N10516, N10318, N6761);
  nand NAND2_3054 (N10518, N10321, N6761);
  nand NAND2_3055 (N10519, N10437, N10325);
  nand NAND2_3056 (N10522, N10438, N10327);
  nand NAND2_3057 (N10525, N10439, N10329);
  nand NAND2_3058 (N10528, N10440, N10331);
  nand NAND2_3059 (N10531, N10441, N10333);
  nand NAND2_3061 (N10535, N10334, N9695);
  nand NAND2_3062 (N10536, N10444, N10338);
  nand NAND2_3063 (N10539, N10445, N10340);
  nand NAND2_3065 (N10543, N10341, N9720);
  nand NAND2_3067 (N10545, N10344, N9726);
  nand NAND2_3074 (N10552, N5856, N10455);
  nand NAND2_3080 (N10558, N10406, N8243);
  nand NAND2_3082 (N10560, N10409, N8244);
  nand NAND2_3084 (N10562, N10412, N8245);
  nand NAND2_3086 (N10564, N10415, N8246);
  nand NAND2_3087 (N10565, N5683, N10465);
  nand NAND2_3089 (N10567, N10419, N8248);
  nand NAND2_3091 (N10569, N10422, N8249);
  nand NAND2_3093 (N10571, N10425, N8250);
  nand NAND2_3095 (N10573, N10428, N8251);
  nand NAND2_3112 (N10609, N5850, N10515);
  nand NAND2_3113 (N10610, N5850, N10517);
  nand NAND2_3114 (N10621, N9149, N10534);
  nand NAND2_3115 (N10626, N9206, N10542);
  nand NAND2_3116 (N10627, N9223, N10544);
  nand NAND2_3120 (N10632, N10552, N10456);
  nand NAND2_3121 (N10637, N5799, N10557);
  nand NAND2_3122 (N10638, N5807, N10559);
  nand NAND2_3123 (N10639, N5821, N10561);
  nand NAND2_3124 (N10640, N5837, N10563);
  nand NAND2_3125 (N10641, N10565, N10466);
  nand NAND2_3126 (N10642, N5632, N10566);
  nand NAND2_3127 (N10643, N5640, N10568);
  nand NAND2_3128 (N10644, N5654, N10570);
  nand NAND2_3129 (N10645, N5670, N10572);
  nand NAND2_3139 (N10672, N10509, N8247);
  nand NAND2_3141 (N10674, N10512, N8247);
  nand NAND2_3142 (N10675, N10609, N10516);
  nand NAND2_3143 (N10678, N10610, N10518);
  nand NAND2_3145 (N10682, N10519, N8242);
  nand NAND2_3147 (N10684, N10522, N8242);
  nand NAND2_3149 (N10686, N10525, N8253);
  nand NAND2_3151 (N10688, N10528, N8253);
  nand NAND2_3153 (N10690, N10531, N9978);
  nand NAND2_3154 (N10691, N10621, N10535);
  nand NAND2_3156 (N10695, N10536, N8252);
  nand NAND2_3158 (N10697, N10539, N8252);
  nand NAND2_3159 (N10698, N10626, N10543);
  nand NAND2_3160 (N10701, N10627, N10545);
  nand NAND2_3168 (N10711, N10637, N10558);
  nand NAND2_3169 (N10712, N10638, N10560);
  nand NAND2_3170 (N10713, N10639, N10562);
  nand NAND2_3171 (N10714, N10640, N10564);
  nand NAND2_3172 (N10715, N10642, N10567);
  nand NAND2_3173 (N10716, N10643, N10569);
  nand NAND2_3174 (N10717, N10644, N10571);
  nand NAND2_3175 (N10718, N10645, N10573);
  nand NAND2_3177 (N10720, N10381, N9244);
  nand NAND2_3181 (N10737, N5683, N10671);
  nand NAND2_3182 (N10738, N5683, N10673);
  nand NAND2_3184 (N10746, N5856, N10681);
  nand NAND2_3185 (N10747, N5856, N10683);
  nand NAND2_3186 (N10748, N6923, N10685);
  nand NAND2_3187 (N10749, N6923, N10687);
  nand NAND2_3188 (N10750, N9685, N10689);
  nand NAND2_3189 (N10753, N7136, N10694);
  nand NAND2_3190 (N10754, N7136, N10696);
  nand NAND2_3196 (N10764, N7180, N10719);
  nand NAND2_3202 (N10770, N10659, N9245);
  nand NAND2_3204 (N10772, N10662, N9246);
  nand NAND2_3206 (N10774, N10665, N9247);
  nand NAND2_3208 (N10776, N10668, N9248);
  nand NAND2_3212 (N10789, N10737, N10672);
  nand NAND2_3213 (N10792, N10738, N10674);
  nand NAND2_3215 (N10797, N10675, N8323);
  nand NAND2_3217 (N10799, N10678, N8323);
  nand NAND2_3218 (N10800, N10746, N10682);
  nand NAND2_3219 (N10803, N10747, N10684);
  nand NAND2_3220 (N10806, N10748, N10686);
  nand NAND2_3221 (N10809, N10749, N10688);
  nand NAND2_3222 (N10812, N10750, N10690);
  nand NAND2_3224 (N10816, N10691, N9741);
  nand NAND2_3225 (N10817, N10753, N10695);
  nand NAND2_3226 (N10820, N10754, N10697);
  nand NAND2_3228 (N10824, N10698, N9244);
  nand NAND2_3230 (N10826, N10701, N9244);
  nand NAND2_3231 (N10827, N10764, N10720);
  nand NAND2_3232 (N10832, N7142, N10769);
  nand NAND2_3233 (N10833, N7149, N10771);
  nand NAND2_3234 (N10834, N7159, N10773);
  nand NAND2_3235 (N10835, N7170, N10775);
  nand NAND2_3241 (N10845, N5789, N10796);
  nand NAND2_3242 (N10846, N5789, N10798);
  nand NAND2_3243 (N10857, N8326, N10815);
  nand NAND2_3244 (N10862, N7180, N10823);
  nand NAND2_3245 (N10863, N7180, N10825);
  nand NAND2_3250 (N10868, N10832, N10770);
  nand NAND2_3251 (N10869, N10833, N10772);
  nand NAND2_3252 (N10870, N10834, N10774);
  nand NAND2_3253 (N10871, N10835, N10776);
  nand NAND2_3255 (N10873, N10789, N8251);
  nand NAND2_3257 (N10875, N10792, N8251);
  nand NAND2_3258 (N10876, N10845, N10797);
  nand NAND2_3259 (N10879, N10846, N10799);
  nand NAND2_3261 (N10883, N10800, N8246);
  nand NAND2_3263 (N10885, N10803, N8246);
  nand NAND2_3265 (N10887, N10806, N9298);
  nand NAND2_3267 (N10889, N10809, N9298);
  nand NAND2_3269 (N10891, N10812, N9741);
  nand NAND2_3270 (N10892, N10857, N10816);
  nand NAND2_3272 (N10896, N10817, N9360);
  nand NAND2_3274 (N10898, N10820, N9360);
  nand NAND2_3275 (N10899, N10862, N10824);
  nand NAND2_3276 (N10902, N10863, N10826);
  nand NAND2_3281 (N10909, N5670, N10872);
  nand NAND2_3282 (N10910, N5670, N10874);
  nand NAND2_3283 (N10915, N5837, N10882);
  nand NAND2_3284 (N10916, N5837, N10884);
  nand NAND2_3285 (N10917, N6912, N10886);
  nand NAND2_3286 (N10918, N6912, N10888);
  nand NAND2_3287 (N10919, N8326, N10890);
  nand NAND2_3288 (N10922, N7125, N10895);
  nand NAND2_3289 (N10923, N7125, N10897);
  nand NAND2_3290 (N10928, N10909, N10873);
  nand NAND2_3291 (N10931, N10910, N10875);
  nand NAND2_3293 (N10935, N10876, N8315);
  nand NAND2_3295 (N10937, N10879, N8315);
  nand NAND2_3296 (N10938, N10915, N10883);
  nand NAND2_3297 (N10941, N10916, N10885);
  nand NAND2_3298 (N10944, N10917, N10887);
  nand NAND2_3299 (N10947, N10918, N10889);
  nand NAND2_3300 (N10950, N10919, N10891);
  nand NAND2_3302 (N10954, N10892, N9252);
  nand NAND2_3303 (N10955, N10922, N10896);
  nand NAND2_3304 (N10958, N10923, N10898);
  nand NAND2_3306 (N10962, N10899, N9248);
  nand NAND2_3308 (N10964, N10902, N9248);
  nand NAND2_3309 (N10969, N5771, N10934);
  nand NAND2_3310 (N10970, N5771, N10936);
  nand NAND2_3311 (N10981, N6957, N10953);
  nand NAND2_3312 (N10986, N7170, N10961);
  nand NAND2_3313 (N10987, N7170, N10963);
  nand NAND2_3315 (N10989, N10928, N8248);
  nand NAND2_3317 (N10991, N10931, N8248);
  nand NAND2_3318 (N10992, N10969, N10935);
  nand NAND2_3319 (N10995, N10970, N10937);
  nand NAND2_3321 (N10999, N10938, N8243);
  nand NAND2_3323 (N11001, N10941, N8243);
  nand NAND2_3325 (N11003, N10944, N9290);
  nand NAND2_3327 (N11005, N10947, N9290);
  nand NAND2_3329 (N11007, N10950, N9252);
  nand NAND2_3330 (N11008, N10981, N10954);
  nand NAND2_3332 (N11012, N10955, N9352);
  nand NAND2_3334 (N11014, N10958, N9352);
  nand NAND2_3335 (N11015, N10986, N10962);
  nand NAND2_3336 (N11018, N10987, N10964);
  nand NAND2_3337 (N11023, N5632, N10988);
  nand NAND2_3338 (N11024, N5632, N10990);
  nand NAND2_3339 (N11027, N5799, N10998);
  nand NAND2_3340 (N11028, N5799, N11000);
  nand NAND2_3341 (N11029, N6894, N11002);
  nand NAND2_3342 (N11030, N6894, N11004);
  nand NAND2_3343 (N11031, N6957, N11006);
  nand NAND2_3344 (N11034, N7107, N11011);
  nand NAND2_3345 (N11035, N7107, N11013);
  nand NAND2_3347 (N11041, N10992, N8294);
  nand NAND2_3349 (N11043, N10995, N8294);
  nand NAND2_3350 (N11044, N11023, N10989);
  nand NAND2_3351 (N11047, N11024, N10991);
  nand NAND2_3352 (N11050, N11027, N10999);
  nand NAND2_3353 (N11053, N11028, N11001);
  nand NAND2_3354 (N11056, N11029, N11003);
  nand NAND2_3355 (N11059, N11030, N11005);
  nand NAND2_3356 (N11062, N11031, N11007);
  nand NAND2_3358 (N11066, N11008, N9249);
  nand NAND2_3359 (N11067, N11034, N11012);
  nand NAND2_3360 (N11070, N11035, N11014);
  nand NAND2_3362 (N11074, N11015, N9245);
  nand NAND2_3364 (N11076, N11018, N9245);
  nand NAND2_3365 (N11077, N5778, N11040);
  nand NAND2_3366 (N11078, N5778, N11042);
  nand NAND2_3367 (N11095, N6929, N11065);
  nand NAND2_3368 (N11098, N7142, N11073);
  nand NAND2_3369 (N11099, N7142, N11075);
  nand NAND2_3370 (N11100, N11077, N11041);
  nand NAND2_3371 (N11103, N11078, N11043);
  nand NAND2_3373 (N11107, N11056, N9294);
  nand NAND2_3375 (N11109, N11059, N9294);
  nand NAND2_3377 (N11111, N11067, N9356);
  nand NAND2_3379 (N11113, N11070, N9356);
  nand NAND2_3381 (N11115, N11044, N8250);
  nand NAND2_3383 (N11117, N11047, N8250);
  nand NAND2_3385 (N11119, N11050, N8245);
  nand NAND2_3387 (N11121, N11053, N8245);
  nand NAND2_3389 (N11123, N11062, N9249);
  nand NAND2_3390 (N11124, N11095, N11066);
  nand NAND2_3391 (N11127, N11098, N11074);
  nand NAND2_3392 (N11130, N11099, N11076);
  nand NAND2_3393 (N11137, N6901, N11106);
  nand NAND2_3394 (N11138, N6901, N11108);
  nand NAND2_3395 (N11139, N7114, N11110);
  nand NAND2_3396 (N11140, N7114, N11112);
  nand NAND2_3397 (N11141, N5654, N11114);
  nand NAND2_3398 (N11142, N5654, N11116);
  nand NAND2_3399 (N11143, N5821, N11118);
  nand NAND2_3400 (N11144, N5821, N11120);
  nand NAND2_3401 (N11145, N6929, N11122);
  nand NAND2_3406 (N11156, N11137, N11107);
  nand NAND2_3407 (N11159, N11138, N11109);
  nand NAND2_3408 (N11162, N11139, N11111);
  nand NAND2_3409 (N11165, N11140, N11113);
  nand NAND2_3410 (N11168, N11141, N11115);
  nand NAND2_3411 (N11171, N11142, N11117);
  nand NAND2_3412 (N11174, N11143, N11119);
  nand NAND2_3413 (N11177, N11144, N11121);
  nand NAND2_3414 (N11180, N11145, N11123);
  nand NAND2_3416 (N11184, N11124, N9251);
  nand NAND2_3418 (N11186, N11127, N9247);
  nand NAND2_3420 (N11188, N11130, N9247);
  nand NAND2_3422 (N11210, N6946, N11183);
  nand NAND2_3423 (N11211, N7159, N11185);
  nand NAND2_3424 (N11212, N7159, N11187);
  nand NAND2_3426 (N11214, N11168, N8249);
  nand NAND2_3428 (N11216, N11171, N8249);
  nand NAND2_3430 (N11218, N11174, N8244);
  nand NAND2_3432 (N11220, N11177, N8244);
  nand NAND2_3442 (N11232, N11180, N9251);
  nand NAND2_3443 (N11233, N11210, N11184);
  nand NAND2_3444 (N11236, N11211, N11186);
  nand NAND2_3445 (N11239, N11212, N11188);
  nand NAND2_3446 (N11242, N5640, N11213);
  nand NAND2_3447 (N11243, N5640, N11215);
  nand NAND2_3448 (N11244, N5807, N11217);
  nand NAND2_3449 (N11245, N5807, N11219);
  nand NAND2_3451 (N11250, N6946, N11231);
  nand NAND2_3454 (N11260, N11242, N11214);
  nand NAND2_3455 (N11261, N11243, N11216);
  nand NAND2_3456 (N11262, N11244, N11218);
  nand NAND2_3457 (N11263, N11245, N11220);
  nand NAND2_3459 (N11265, N11233, N9250);
  nand NAND2_3461 (N11268, N11236, N9246);
  nand NAND2_3463 (N11270, N11239, N9246);
  nand NAND2_3464 (N11272, N11250, N11232);
  nand NAND2_3469 (N11282, N6936, N11264);
  nand NAND2_3471 (N11284, N7149, N11267);
  nand NAND2_3472 (N11285, N7149, N11269);
  nand NAND2_3477 (N11291, N11272, N9250);
  nand NAND2_3478 (N11292, N11282, N11265);
  nand NAND2_3479 (N11293, N11284, N11268);
  nand NAND2_3480 (N11294, N11285, N11270);
  nand NAND2_3481 (N11295, N6936, N11290);
  nand NAND2_3487 (N11307, N11295, N11291);
  nand NAND2_3490 (N11312, N11302, N11246);
  nand NAND2_3491 (N11313, N11299, N10836);
  nand NAND2_3496 (N11320, N11205, N11315);
  nand NAND2_3497 (N11321, N10739, N11314);
  nand NAND2_3499 (N11327, N11312, N11320);
  nand NAND2_3500 (N11328, N11313, N11321);
  nand NAND2_3501 (N11329, N11317, N11286);
  nand NAND2_3505 (N11335, N11257, N11331);
  nand NAND2_3506 (N11336, N11323, N11283);
  nand NAND2_3508 (N11338, N11329, N11335);
  nand NAND2_3509 (N11339, N11252, N11337);
  nand NAND2_3511 (N11341, N11336, N11339);
  nor NOR2_230 (N1708, N957, N38);
  nor NOR2_784 (N3507, N1167, N2866);
  nor NOR2_786 (N3515, N644, N2619);
  nor NOR2_824 (N3625, N734, N2488);
  nor NOR2_825 (N3628, N708, N2554);
  nor NOR2_1161 (N4844, N3273, N786);
  nor NOR2_1193 (N4940, N3390, N845);
  nor NOR2_1223 (N5030, N814, N3315);
  nor NOR2_1610 (N6217, N2674, N4769);
  nor NOR2_2045 (N8208, N3173, N6844);
  nor NOR2_2421 (N9111, N4549, N8345);
  nor NOR2_2431 (N9173, N4661, N8441);
  nor NOR2_2458 (N9256, N8861, N8280);
  nor NOR2_2459 (N9257, N8862, N8281);
  nor NOR2_2460 (N9258, N8863, N8282);
  nor NOR2_2461 (N9259, N8864, N8283);
  nor NOR2_2462 (N9260, N8865, N8284);
  nor NOR2_2463 (N9261, N8866, N8285);
  nor NOR2_2513 (N9367, N8991, N8483);
  nor NOR2_2514 (N9368, N8992, N8484);
  nor NOR2_2533 (N9400, N9024, N8539);
  nor NOR2_2534 (N9401, N9025, N8540);
  nor NOR2_2543 (N9417, N9053, N8578);
  nor NOR2_2544 (N9418, N9054, N8579);
  nor NOR2_2724 (N9800, N9602, N9369);
  nor NOR2_2725 (N9801, N9603, N9370);
  nor NOR2_2726 (N9802, N9604, N9371);
  nor NOR2_2727 (N9803, N9605, N9372);
  nor NOR2_2731 (N9813, N9612, N9396);
  nor NOR2_2732 (N9814, N9613, N9397);
  nor NOR2_2733 (N9815, N9614, N9398);
  nor NOR2_2734 (N9816, N9615, N9399);
  nor NOR2_2739 (N9827, N9621, N9419);
  nor NOR2_2740 (N9828, N9622, N9420);
  nor NOR2_2741 (N9829, N9623, N9421);
  nor NOR2_2742 (N9830, N9624, N9422);
  nor NOR3_2032 (N8131, N3101, N6777, N6778);
  nor NOR3_2037 (N8156, N3169, N6839, N6840);
  nor NOR3_2040 (N8183, N3189, N6859, N6860);
  nor NOR3_2419 (N9103, N4545, N8340, N8341);
  nor NOR3_2424 (N9146, N4566, N8355, N8356);
  nor NOR3_2429 (N9165, N4657, N8436, N8437);
  nor NOR3_2440 (N9220, N4678, N8454, N8455);
  nor NOR4_2033 (N8134, N3097, N6770, N6771, N6772);
  nor NOR4_2041 (N8186, N3185, N6852, N6853, N6854);
  nor NOR4_2425 (N9149, N4563, N8352, N8353, N8354);
  nor NOR4_2441 (N9223, N4675, N8451, N8452, N8453);
  not NOT1_3 (N467, N57);
  not NOT1_43 (N582, N15);
  not NOT1_44 (N585, N5);
  not NOT1_48 (N599, N289);
  not NOT1_49 (N604, N299);
  not NOT1_50 (N609, N303);
  not NOT1_56 (N641, N245);
  not NOT1_57 (N642, N248);
  not NOT1_59 (N644, N251);
  not NOT1_60 (N651, N254);
  not NOT1_62 (N660, N257);
  not NOT1_63 (N666, N260);
  not NOT1_64 (N672, N263);
  not NOT1_65 (N673, N267);
  not NOT1_66 (N674, N106);
  not NOT1_71 (N695, N18);
  not NOT1_73 (N705, N271);
  not NOT1_74 (N706, N274);
  not NOT1_76 (N708, N277);
  not NOT1_77 (N715, N280);
  not NOT1_78 (N721, N283);
  not NOT1_79 (N727, N286);
  not NOT1_81 (N734, N293);
  not NOT1_82 (N742, N296);
  not NOT1_86 (N758, N307);
  not NOT1_87 (N759, N310);
  not NOT1_88 (N762, N313);
  not NOT1_89 (N768, N316);
  not NOT1_90 (N774, N319);
  not NOT1_91 (N780, N322);
  not NOT1_92 (N786, N325);
  not NOT1_93 (N794, N328);
  not NOT1_94 (N800, N331);
  not NOT1_95 (N806, N334);
  not NOT1_96 (N812, N337);
  not NOT1_98 (N814, N340);
  not NOT1_99 (N821, N343);
  not NOT1_100 (N827, N346);
  not NOT1_101 (N833, N349);
  not NOT1_102 (N839, N352);
  not NOT1_103 (N845, N355);
  not NOT1_104 (N853, N358);
  not NOT1_105 (N859, N361);
  not NOT1_106 (N865, N364);
  not NOT1_109 (N882, N528);
  not NOT1_110 (N883, N578);
  not NOT1_111 (N884, N575);
  not NOT1_112 (N885, N494);
  not NOT1_117 (N957, N688);
  not NOT1_126 (N1115, N367);
  not NOT1_146 (N1222, N1028);
  not NOT1_224 (N1113, N1109);
  not NOT1_256 (N1821, N700);
  not NOT1_257 (N1822, N38);
  not NOT1_401 (N2117, N1708);
  not NOT1_402 (N2171, N1029);
  not NOT1_560 (N2537, N1537);
  not NOT1_674 (N3073, N628);
  not NOT1_675 (N3080, N2441);
  not NOT1_686 (N3135, N2523);
  not NOT1_694 (N3167, N2778);
  not NOT1_751 (N3380, N2781);
  not NOT1_767 (N3452, N2790);
  not NOT1_768 (N3453, N2793);
  not NOT1_777 (N3486, N2796);
  not NOT1_797 (N3551, N2766);
  not NOT1_798 (N3552, N2769);
  not NOT1_804 (N3569, N2772);
  not NOT1_805 (N3570, N2775);
  not NOT1_876 (N3781, N2784);
  not NOT1_877 (N3782, N2787);
  not NOT1_916 (N3954, N2257);
  not NOT1_932 (N4464, N2644);
  not NOT1_934 (N4466, N2638);
  not NOT1_936 (N4468, N2632);
  not NOT1_938 (N4470, N2626);
  not NOT1_940 (N4472, N2619);
  not NOT1_941 (N4473, N3122);
  not NOT1_965 (N4497, N2450);
  not NOT1_966 (N4498, N2446);
  not NOT1_967 (N4499, N2458);
  not NOT1_968 (N4500, N2454);
  not NOT1_969 (N4501, N2554);
  not NOT1_971 (N4503, N2567);
  not NOT1_972 (N4504, N2561);
  not NOT1_973 (N4505, N2482);
  not NOT1_974 (N4506, N2573);
  not NOT1_976 (N4508, N2508);
  not NOT1_978 (N4510, N2502);
  not NOT1_980 (N4512, N2496);
  not NOT1_990 (N4522, N2488);
  not NOT1_1011 (N4543, N3625);
  not NOT1_1020 (N4575, N2674);
  not NOT1_1030 (N4611, N2761);
  not NOT1_1031 (N4612, N2478);
  not NOT1_1032 (N4613, N2757);
  not NOT1_1033 (N4614, N2474);
  not NOT1_1034 (N4615, N2753);
  not NOT1_1035 (N4616, N2470);
  not NOT1_1036 (N4617, N2745);
  not NOT1_1037 (N4618, N2462);
  not NOT1_1038 (N4619, N2741);
  not NOT1_1039 (N4620, N2550);
  not NOT1_1040 (N4621, N2737);
  not NOT1_1041 (N4622, N2546);
  not NOT1_1042 (N4623, N2733);
  not NOT1_1043 (N4624, N2542);
  not NOT1_1044 (N4625, N2749);
  not NOT1_1045 (N4626, N2466);
  not NOT1_1046 (N4627, N2729);
  not NOT1_1047 (N4628, N2538);
  not NOT1_1048 (N4629, N2704);
  not NOT1_1050 (N4631, N2700);
  not NOT1_1052 (N4633, N2696);
  not NOT1_1055 (N4636, N2688);
  not NOT1_1061 (N4642, N2692);
  not NOT1_1062 (N4643, N2670);
  not NOT1_1064 (N4645, N2666);
  not NOT1_1066 (N4647, N2662);
  not NOT1_1068 (N4649, N2658);
  not NOT1_1070 (N4651, N2654);
  not NOT1_1072 (N4653, N3375);
  not NOT1_1088 (N4699, N3783);
  not NOT1_1089 (N4700, N3786);
  not NOT1_1099 (N4743, N3789);
  not NOT1_1101 (N4745, N2604);
  not NOT1_1103 (N4747, N2611);
  not NOT1_1104 (N4748, N2607);
  not NOT1_1105 (N4749, N2615);
  not NOT1_1124 (N4768, N2680);
  not NOT1_1132 (N4781, N3885);
  not NOT1_1133 (N4782, N3888);
  not NOT1_1134 (N4783, N3891);
  not NOT1_1138 (N3126, N3507);
  not NOT1_1140 (N4795, N3515);
  not NOT1_1150 (N4813, N3628);
  not NOT1_1351 (N5324, N4193);
  not NOT1_1372 (N5469, N4303);
  not NOT1_1400 (N5735, N5177);
  not NOT1_1410 (N5769, N4803);
  not NOT1_1411 (N5770, N4806);
  not NOT1_1430 (N5943, N3178);
  not NOT1_1432 (N5945, N3293);
  not NOT1_1434 (N5947, N3287);
  not NOT1_1436 (N5949, N3281);
  not NOT1_1438 (N5951, N3273);
  not NOT1_1440 (N5953, N3267);
  not NOT1_1442 (N5955, N3355);
  not NOT1_1444 (N5957, N3349);
  not NOT1_1446 (N5959, N3343);
  not NOT1_1448 (N5966, N4844);
  not NOT1_1475 (N6023, N3448);
  not NOT1_1477 (N6025, N3444);
  not NOT1_1479 (N6027, N3440);
  not NOT1_1481 (N6029, N3432);
  not NOT1_1483 (N6031, N3428);
  not NOT1_1484 (N6032, N3311);
  not NOT1_1485 (N6033, N3424);
  not NOT1_1486 (N6034, N3307);
  not NOT1_1487 (N6035, N3420);
  not NOT1_1488 (N6036, N3303);
  not NOT1_1489 (N6037, N3436);
  not NOT1_1491 (N6039, N3416);
  not NOT1_1492 (N6040, N3299);
  not NOT1_1499 (N6061, N3410);
  not NOT1_1501 (N6063, N3404);
  not NOT1_1503 (N6065, N3398);
  not NOT1_1505 (N6067, N3390);
  not NOT1_1507 (N6069, N3384);
  not NOT1_1509 (N6071, N3334);
  not NOT1_1511 (N6073, N3328);
  not NOT1_1513 (N6075, N3322);
  not NOT1_1515 (N6077, N3315);
  not NOT1_1516 (N6078, N4940);
  not NOT1_1526 (N6096, N3340);
  not NOT1_1532 (N6102, N4997);
  not NOT1_1559 (N6135, N3247);
  not NOT1_1564 (N6148, N3482);
  not NOT1_1565 (N6149, N3263);
  not NOT1_1566 (N6150, N3478);
  not NOT1_1567 (N6151, N3259);
  not NOT1_1568 (N6152, N3474);
  not NOT1_1569 (N6153, N3255);
  not NOT1_1570 (N6154, N3466);
  not NOT1_1572 (N6156, N3462);
  not NOT1_1574 (N6158, N3458);
  not NOT1_1576 (N6160, N3454);
  not NOT1_1578 (N6162, N3470);
  not NOT1_1579 (N6163, N3251);
  not NOT1_1581 (N6165, N3381);
  not NOT1_1596 (N6191, N4784);
  not NOT1_1600 (N6195, N3114);
  not NOT1_1604 (N6203, N3202);
  not NOT1_1622 (N6235, N5030);
  not NOT1_1749 (N6761, N5850);
  not NOT1_1780 (N6797, N5736);
  not NOT1_1781 (N6800, N5740);
  not NOT1_1782 (N6803, N5747);
  not NOT1_1783 (N6806, N5751);
  not NOT1_1784 (N6809, N5758);
  not NOT1_1785 (N6812, N5762);
  not NOT1_1854 (N6968, N4769);
  not NOT1_1855 (N6969, N4555);
  not NOT1_1898 (N7187, N4667);
  not NOT1_1899 (N7188, N6079);
  not NOT1_1900 (N7191, N6083);
  not NOT1_1921 (N7325, N6127);
  not NOT1_1922 (N7328, N6131);
  not NOT1_1924 (N7334, N6137);
  not NOT1_1925 (N7337, N6141);
  not NOT1_1937 (N7378, N6166);
  not NOT1_1938 (N7381, N6170);
  not NOT1_1939 (N7384, N6177);
  not NOT1_1969 (N7477, N6196);
  not NOT1_1970 (N7478, N6199);
  not NOT1_1996 (N7552, N6217);
  not NOT1_1998 (N7556, N6249);
  not NOT1_1999 (N7557, N6252);
  not NOT1_2000 (N7558, N6243);
  not NOT1_2001 (N7559, N6246);
  not NOT1_2007 (N7573, N4687);
  not NOT1_2010 (N7580, N6263);
  not NOT1_2011 (N7581, N6266);
  not NOT1_2052 (N8242, N5856);
  not NOT1_2053 (N8243, N5799);
  not NOT1_2054 (N8244, N5807);
  not NOT1_2055 (N8245, N5821);
  not NOT1_2056 (N8246, N5837);
  not NOT1_2057 (N8247, N5683);
  not NOT1_2058 (N8248, N5632);
  not NOT1_2059 (N8249, N5640);
  not NOT1_2060 (N8250, N5654);
  not NOT1_2061 (N8251, N5670);
  not NOT1_2062 (N8252, N7136);
  not NOT1_2063 (N8253, N6923);
  not NOT1_2064 (N8254, N6762);
  not NOT1_2069 (N8274, N5744);
  not NOT1_2071 (N8276, N5755);
  not NOT1_2073 (N8278, N5766);
  not NOT1_2081 (N8288, N6845);
  not NOT1_2082 (N8294, N5778);
  not NOT1_2088 (N8315, N5771);
  not NOT1_2093 (N8323, N5789);
  not NOT1_2181 (N8457, N7194);
  not NOT1_2182 (N8460, N7198);
  not NOT1_2183 (N8463, N7205);
  not NOT1_2184 (N8466, N7209);
  not NOT1_2185 (N8469, N6087);
  not NOT1_2223 (N8519, N7314);
  not NOT1_2224 (N8522, N7318);
  not NOT1_2229 (N8537, N6145);
  not NOT1_2242 (N8555, N7387);
  not NOT1_2243 (N8558, N7394);
  not NOT1_2244 (N8561, N7398);
  not NOT1_2245 (N8564, N6174);
  not NOT1_2262 (N8607, N7441);
  not NOT1_2264 (N8609, N7444);
  not NOT1_2308 (N8717, N5960);
  not NOT1_2314 (N8733, N7574);
  not NOT1_2315 (N8734, N7577);
  not NOT1_2322 (N8753, N7560);
  not NOT1_2323 (N8754, N7563);
  not NOT1_2324 (N8755, N7566);
  not NOT1_2325 (N8756, N7569);
  not NOT1_2345 (N8814, N7588);
  not NOT1_2346 (N8815, N7591);
  not NOT1_2347 (N8816, N7582);
  not NOT1_2348 (N8817, N7585);
  not NOT1_2351 (N8857, N7609);
  not NOT1_2358 (N8871, N7655);
  not NOT1_2361 (N8879, N8146);
  not NOT1_2363 (N8881, N8156);
  not NOT1_2365 (N8883, N8204);
  not NOT1_2367 (N7650, N8208);
  not NOT1_2380 (N8959, N7852);
  not NOT1_2398 (N9066, N8114);
  not NOT1_2401 (N9071, N8117);
  not NOT1_2402 (N9072, N8131);
  not NOT1_2404 (N9074, N7613);
  not NOT1_2405 (N9077, N8134);
  not NOT1_2410 (N9087, N8166);
  not NOT1_2413 (N9092, N8169);
  not NOT1_2414 (N9093, N8183);
  not NOT1_2416 (N9095, N7659);
  not NOT1_2417 (N9098, N8186);
  not NOT1_2449 (N9244, N7180);
  not NOT1_2450 (N9245, N7142);
  not NOT1_2451 (N9246, N7149);
  not NOT1_2452 (N9247, N7159);
  not NOT1_2453 (N9248, N7170);
  not NOT1_2454 (N9249, N6929);
  not NOT1_2455 (N9250, N6936);
  not NOT1_2456 (N9251, N6946);
  not NOT1_2457 (N9252, N6957);
  not NOT1_2464 (N9262, N8627);
  not NOT1_2472 (N9276, N8333);
  not NOT1_2478 (N9290, N6894);
  not NOT1_2480 (N9294, N6901);
  not NOT1_2483 (N9298, N6912);
  not NOT1_2495 (N9323, N8727);
  not NOT1_2496 (N9324, N8730);
  not NOT1_2497 (N9326, N8405);
  not NOT1_2501 (N9352, N7107);
  not NOT1_2503 (N9356, N7114);
  not NOT1_2506 (N9360, N7125);
  not NOT1_2509 (N9363, N7202);
  not NOT1_2511 (N9365, N7213);
  not NOT1_2519 (N9375, N8497);
  not NOT1_2525 (N9392, N7322);
  not NOT1_2527 (N9394, N7331);
  not NOT1_2535 (N9402, N8541);
  not NOT1_2538 (N9412, N8811);
  not NOT1_2539 (N9413, N7391);
  not NOT1_2541 (N9415, N7402);
  not NOT1_2593 (N9541, N9275);
  not NOT1_2598 (N9557, N8898);
  not NOT1_2600 (N9561, N9099);
  not NOT1_2602 (N9563, N9103);
  not NOT1_2604 (N9565, N9107);
  not NOT1_2606 (N8924, N9111);
  not NOT1_2611 (N9575, N8902);
  not NOT1_2613 (N9581, N8950);
  not NOT1_2614 (N9582, N8956);
  not NOT1_2617 (N9592, N9161);
  not NOT1_2619 (N9594, N9165);
  not NOT1_2621 (N9596, N9169);
  not NOT1_2623 (N8996, N9173);
  not NOT1_2631 (N9608, N8966);
  not NOT1_2637 (N9616, N9029);
  not NOT1_2638 (N9617, N9035);
  not NOT1_2649 (N9645, N9068);
  not NOT1_2655 (N9659, N9079);
  not NOT1_2660 (N9666, N9089);
  not NOT1_2670 (N9690, N9146);
  not NOT1_2672 (N9692, N8931);
  not NOT1_2673 (N9695, N9149);
  not NOT1_2680 (N9715, N9203);
  not NOT1_2683 (N9720, N9206);
  not NOT1_2684 (N9721, N9220);
  not NOT1_2686 (N9723, N9005);
  not NOT1_2687 (N9726, N9223);
  not NOT1_2694 (N9737, N9555);
  not NOT1_2695 (N9738, N9556);
  not NOT1_2698 (N9741, N8326);
  not NOT1_2709 (N9769, N9307);
  not NOT1_2714 (N9784, N9478);
  not NOT1_2728 (N9805, N9485);
  not NOT1_2729 (N9806, N9488);
  not NOT1_2737 (N9825, N9517);
  not NOT1_2738 (N9826, N9520);
  not NOT1_2743 (N9835, N9426);
  not NOT1_2745 (N9837, N9429);
  not NOT1_2756 (N9892, N9799);
  not NOT1_2760 (N9896, N9766);
  not NOT1_2761 (N9897, N9626);
  not NOT1_2763 (N9899, N9629);
  not NOT1_2765 (N9901, N9632);
  not NOT1_2767 (N9903, N9635);
  not NOT1_2769 (N9905, N9543);
  not NOT1_2770 (N9906, N9650);
  not NOT1_2772 (N9908, N9653);
  not NOT1_2774 (N9910, N9656);
  not NOT1_2776 (N9917, N9551);
  not NOT1_2782 (N9938, N9698);
  not NOT1_2786 (N9947, N9702);
  not NOT1_2789 (N9953, N9727);
  not NOT1_2793 (N9957, N9642);
  not NOT1_2795 (N9959, N9646);
  not NOT1_2799 (N9967, N9663);
  not NOT1_2801 (N9969, N9667);
  not NOT1_2803 (N9971, N9671);
  not NOT1_2807 (N9975, N9679);
  not NOT1_2809 (N9977, N9682);
  not NOT1_2810 (N9978, N9685);
  not NOT1_2817 (N9995, N9707);
  not NOT1_2822 (N10002, N9717);
  not NOT1_2837 (N10023, N9945);
  not NOT1_2838 (N10024, N9946);
  not NOT1_2840 (N10026, N9923);
  not NOT1_2841 (N10028, N9924);
  not NOT1_2855 (N10053, N9817);
  not NOT1_2894 (N10124, N9925);
  not NOT1_2896 (N10131, N9932);
  not NOT1_2897 (N10132, N9935);
  not NOT1_2900 (N10135, N9983);
  not NOT1_2902 (N10137, N9986);
  not NOT1_2909 (N10156, N9989);
  not NOT1_2911 (N10158, N9992);
  not NOT1_2913 (N10160, N9949);
  not NOT1_2915 (N10162, N10007);
  not NOT1_2917 (N10164, N10010);
  not NOT1_2921 (N10176, N9961);
  not NOT1_2923 (N10178, N9964);
  not NOT1_2930 (N10195, N9979);
  not NOT1_2934 (N10203, N9999);
  not NOT1_2936 (N10205, N10003);
  not NOT1_2949 (N10241, N10070);
  not NOT1_2950 (N10242, N10073);
  not NOT1_2969 (N10283, N10119);
  not NOT1_2987 (N10314, N10170);
  not NOT1_2989 (N10316, N10173);
  not NOT1_2993 (N10324, N10180);
  not NOT1_2995 (N10326, N10183);
  not NOT1_2997 (N10328, N10186);
  not NOT1_2999 (N10330, N10189);
  not NOT1_3001 (N10332, N10192);
  not NOT1_3004 (N10337, N10197);
  not NOT1_3006 (N10339, N10200);
  not NOT1_3041 (N10450, N10296);
  not NOT1_3043 (N10455, N10148);
  not NOT1_3045 (N10465, N10141);
  not NOT1_3047 (N10479, N10116);
  not NOT1_3048 (N10497, N10301);
  not NOT1_3051 (N10515, N10318);
  not NOT1_3053 (N10517, N10321);
  not NOT1_3060 (N10534, N10334);
  not NOT1_3064 (N10542, N10341);
  not NOT1_3066 (N10544, N10344);
  not NOT1_3069 (N10547, N10391);
  not NOT1_3072 (N10550, N10354);
  not NOT1_3079 (N10557, N10406);
  not NOT1_3081 (N10559, N10409);
  not NOT1_3083 (N10561, N10412);
  not NOT1_3085 (N10563, N10415);
  not NOT1_3088 (N10566, N10419);
  not NOT1_3090 (N10568, N10422);
  not NOT1_3092 (N10570, N10425);
  not NOT1_3094 (N10572, N10428);
  not NOT1_3096 (N10574, N10399);
  not NOT1_3097 (N10575, N10402);
  not NOT1_3098 (N10576, N10388);
  not NOT1_3102 (N10583, N10367);
  not NOT1_3105 (N10589, N10375);
  not NOT1_3138 (N10671, N10509);
  not NOT1_3140 (N10673, N10512);
  not NOT1_3144 (N10681, N10519);
  not NOT1_3146 (N10683, N10522);
  not NOT1_3148 (N10685, N10525);
  not NOT1_3150 (N10687, N10528);
  not NOT1_3152 (N10689, N10531);
  not NOT1_3155 (N10694, N10536);
  not NOT1_3157 (N10696, N10539);
  not NOT1_3176 (N10719, N10381);
  not NOT1_3178 (N10729, N10647);
  not NOT1_3201 (N10769, N10659);
  not NOT1_3203 (N10771, N10662);
  not NOT1_3205 (N10773, N10665);
  not NOT1_3207 (N10775, N10668);
  not NOT1_3211 (N10784, N10652);
  not NOT1_3214 (N10796, N10675);
  not NOT1_3216 (N10798, N10678);
  not NOT1_3223 (N10815, N10691);
  not NOT1_3227 (N10823, N10698);
  not NOT1_3229 (N10825, N10701);
  not NOT1_3236 (N10836, N10739);
  not NOT1_3254 (N10872, N10789);
  not NOT1_3256 (N10874, N10792);
  not NOT1_3260 (N10882, N10800);
  not NOT1_3262 (N10884, N10803);
  not NOT1_3264 (N10886, N10806);
  not NOT1_3266 (N10888, N10809);
  not NOT1_3268 (N10890, N10812);
  not NOT1_3271 (N10895, N10817);
  not NOT1_3273 (N10897, N10820);
  not NOT1_3292 (N10934, N10876);
  not NOT1_3294 (N10936, N10879);
  not NOT1_3301 (N10953, N10892);
  not NOT1_3305 (N10961, N10899);
  not NOT1_3307 (N10963, N10902);
  not NOT1_3314 (N10988, N10928);
  not NOT1_3316 (N10990, N10931);
  not NOT1_3320 (N10998, N10938);
  not NOT1_3322 (N11000, N10941);
  not NOT1_3324 (N11002, N10944);
  not NOT1_3326 (N11004, N10947);
  not NOT1_3328 (N11006, N10950);
  not NOT1_3331 (N11011, N10955);
  not NOT1_3333 (N11013, N10958);
  not NOT1_3346 (N11040, N10992);
  not NOT1_3348 (N11042, N10995);
  not NOT1_3357 (N11065, N11008);
  not NOT1_3361 (N11073, N11015);
  not NOT1_3363 (N11075, N11018);
  not NOT1_3372 (N11106, N11056);
  not NOT1_3374 (N11108, N11059);
  not NOT1_3376 (N11110, N11067);
  not NOT1_3378 (N11112, N11070);
  not NOT1_3380 (N11114, N11044);
  not NOT1_3382 (N11116, N11047);
  not NOT1_3384 (N11118, N11050);
  not NOT1_3386 (N11120, N11053);
  not NOT1_3388 (N11122, N11062);
  not NOT1_3415 (N11183, N11124);
  not NOT1_3417 (N11185, N11127);
  not NOT1_3419 (N11187, N11130);
  not NOT1_3425 (N11213, N11168);
  not NOT1_3427 (N11215, N11171);
  not NOT1_3429 (N11217, N11174);
  not NOT1_3431 (N11219, N11177);
  not NOT1_3441 (N11231, N11180);
  not NOT1_3450 (N11246, N11205);
  not NOT1_3458 (N11264, N11233);
  not NOT1_3460 (N11267, N11236);
  not NOT1_3462 (N11269, N11239);
  not NOT1_3465 (N11277, N11261);
  not NOT1_3467 (N11279, N11263);
  not NOT1_3470 (N11283, N11252);
  not NOT1_3473 (N11286, N11257);
  not NOT1_3476 (N11290, N11272);
  not NOT1_3482 (N11296, N11292);
  not NOT1_3483 (N11297, N11294);
  not NOT1_3492 (N11314, N11299);
  not NOT1_3493 (N11315, N11302);
  not NOT1_3502 (N11331, N11317);
  not NOT1_3503 (N11333, N11327);
  not NOT1_3504 (N11334, N11328);
  not NOT1_3507 (N11337, N11323);
  not NOT1_3510 (N11340, N11338);
  not NOT1_3512 (N11342, N11341);
  or OR2_407 (N2239, N695, N1782);
  or OR2_409 (N2241, N695, N1793);
  or OR2_410 (N2242, N695, N1794);
  or OR2_411 (N2243, N695, N1795);
  or OR2_412 (N2244, N695, N1796);
  or OR2_413 (N2245, N695, N1797);
  or OR2_414 (N2246, N695, N1798);
  or OR2_415 (N2247, N695, N1811);
  or OR2_416 (N2248, N695, N1812);
  or OR2_417 (N2249, N695, N1813);
  or OR2_418 (N2250, N695, N1814);
  or OR2_419 (N2251, N695, N1815);
  or OR2_420 (N2252, N695, N1816);
  or OR2_421 (N2253, N695, N1817);
  or OR2_422 (N2254, N695, N1818);
  or OR2_423 (N2255, N695, N1819);
  or OR2_424 (N2256, N695, N1820);
  or OR2_477 (N2348, N695, N1957);
  or OR2_478 (N2349, N695, N1958);
  or OR2_479 (N2350, N695, N1959);
  or OR2_480 (N2351, N695, N1960);
  or OR2_481 (N2352, N695, N1961);
  or OR2_482 (N2353, N695, N1962);
  or OR2_483 (N2354, N695, N1963);
  or OR2_561 (N2538, N2278, N1858);
  or OR2_562 (N2542, N2279, N1859);
  or OR2_563 (N2546, N2280, N1860);
  or OR2_564 (N2550, N2281, N1861);
  or OR2_565 (N2554, N2278, N1863);
  or OR2_566 (N2561, N2279, N1864);
  or OR2_567 (N2567, N2280, N1865);
  or OR2_568 (N2573, N2281, N1866);
  or OR2_569 (N2604, N2338, N1927);
  or OR2_570 (N2607, N2339, N1928);
  or OR2_571 (N2611, N2340, N1929);
  or OR2_572 (N2615, N2341, N1930);
  or OR2_580 (N2654, N2359, N1990);
  or OR2_581 (N2658, N2360, N1991);
  or OR2_582 (N2662, N2361, N1992);
  or OR2_583 (N2666, N2362, N1993);
  or OR2_584 (N2670, N2363, N1994);
  or OR2_585 (N2674, N2366, N18);
  or OR2_586 (N2680, N2367, N18);
  or OR2_587 (N2688, N2374, N2010);
  or OR2_588 (N2692, N2375, N2011);
  or OR2_589 (N2696, N2376, N2012);
  or OR2_590 (N2700, N2377, N2013);
  or OR2_591 (N2704, N2378, N2014);
  or OR2_593 (N2729, N2429, N2065);
  or OR2_594 (N2733, N2430, N2066);
  or OR2_595 (N2737, N2431, N2067);
  or OR2_596 (N2741, N2432, N2068);
  or OR2_597 (N2745, N2433, N2069);
  or OR2_598 (N2749, N2434, N2070);
  or OR2_599 (N2753, N2435, N2071);
  or OR2_600 (N2757, N2436, N2072);
  or OR2_601 (N2761, N2437, N2073);
  or OR2_607 (N2778, N2277, N1862);
  or OR2_608 (N2781, N2358, N1989);
  or OR2_609 (N2784, N2365, N1996);
  or OR2_610 (N2787, N2364, N1995);
  or OR2_611 (N2790, N2337, N1926);
  or OR2_612 (N2793, N2277, N1857);
  or OR2_613 (N2796, N2428, N2064);
  or OR2_713 (N3247, N2913, N2299);
  or OR2_714 (N3251, N2914, N2300);
  or OR2_715 (N3255, N2915, N2301);
  or OR2_716 (N3259, N2916, N2302);
  or OR2_717 (N3263, N2917, N2303);
  or OR2_718 (N3267, N2918, N2299);
  or OR2_719 (N3273, N2919, N2300);
  or OR2_720 (N3281, N2920, N2301);
  or OR2_721 (N3287, N2921, N2302);
  or OR2_722 (N3293, N2922, N2303);
  or OR2_723 (N3299, N2924, N2322);
  or OR2_724 (N3303, N2925, N2323);
  or OR2_725 (N3307, N2926, N2324);
  or OR2_726 (N3311, N2927, N2325);
  or OR2_727 (N3315, N2929, N2322);
  or OR2_728 (N3322, N2930, N2323);
  or OR2_729 (N3328, N2931, N2324);
  or OR2_730 (N3334, N2932, N2325);
  or OR2_731 (N3340, N2934, N1927);
  or OR2_732 (N3343, N2935, N1928);
  or OR2_733 (N3349, N2936, N1929);
  or OR2_734 (N3355, N2937, N1930);
  or OR2_753 (N3384, N3005, N2010);
  or OR2_754 (N3390, N3006, N2011);
  or OR2_755 (N3398, N3007, N2012);
  or OR2_756 (N3404, N3008, N2013);
  or OR2_757 (N3410, N3009, N2014);
  or OR2_758 (N3416, N3021, N2397);
  or OR2_759 (N3420, N3022, N2398);
  or OR2_760 (N3424, N3023, N2399);
  or OR2_761 (N3428, N3024, N2400);
  or OR2_762 (N3432, N3025, N2401);
  or OR2_763 (N3436, N3026, N2402);
  or OR2_764 (N3440, N3027, N2403);
  or OR2_765 (N3444, N3028, N2404);
  or OR2_766 (N3448, N3029, N2405);
  or OR2_769 (N3454, N3034, N2420);
  or OR2_770 (N3458, N3035, N2421);
  or OR2_771 (N3462, N3036, N2422);
  or OR2_772 (N3466, N3037, N2423);
  or OR2_773 (N3470, N3038, N2424);
  or OR2_774 (N3474, N3039, N2425);
  or OR2_775 (N3478, N3040, N2426);
  or OR2_776 (N3482, N3041, N2427);
  or OR2_878 (N3783, N2928, N2321);
  or OR2_879 (N3786, N2933, N1926);
  or OR2_880 (N3789, N2923, N2321);
  or OR2_912 (N3885, N3033, N2367);
  or OR2_913 (N3888, N3032, N2418);
  or OR2_914 (N3891, N3020, N2396);
  or OR2_921 (N4193, N1649, N3379);
  or OR2_1135 (N4784, N3126, N3122);
  or OR2_2017 (N7613, N3107, N6782);
  or OR2_2022 (N7659, N3195, N6864);
  or OR2_2376 (N8931, N4570, N8357);
  or OR2_2377 (N8943, N7825, N8404);
  or OR2_2389 (N9005, N4682, N8456);
  or OR2_2400 (N9068, N7613, N6783);
  or OR2_2406 (N9079, N7650, N6865);
  or OR2_2412 (N9089, N7659, N6866);
  or OR2_2465 (N9265, N7649, N8874);
  or OR2_2647 (N9635, N5960, N9288);
  or OR2_2663 (N9671, N8924, N8346);
  or OR2_2668 (N9682, N8931, N9318);
  or OR2_2676 (N9707, N8996, N8442);
  or OR2_2682 (N9717, N9005, N8518);
  or OR2_2701 (N9758, N8898, N9560);
  or OR2_2716 (N9786, N8950, N9585);
  or OR2_2718 (N9791, N8963, N9591);
  or OR2_2736 (N9820, N9029, N9618);
  or OR2_2779 (N9925, N8902, N9767);
  or OR2_2943 (N10233, N10139, N10054);
  or OR2_2982 (N10301, N10230, N10133);
  or OR2_3010 (N10350, N10266, N10105);
  or OR2_3011 (N10351, N10267, N10106);
  or OR2_3012 (N10352, N10268, N10107);
  or OR2_3013 (N10353, N10269, N10108);
  or OR2_3017 (N10367, N7609, N10282);
  or OR2_3018 (N10375, N7655, N10291);
  or OR2_3019 (N10381, N10292, N10130);
  or OR2_3027 (N10415, N3202, N10290);
  or OR2_3031 (N10428, N3114, N10281);
  or OR2_3117 (N10628, N10546, N10451);
  or OR2_3133 (N10652, N8966, N10598);
  or OR2_3137 (N10668, N4687, N10597);
  or OR2_3161 (N10704, N10629, N10548);
  or OR2_3163 (N10706, N10631, N10551);
  or OR2_3191 (N10759, N10705, N10549);
  or OR2_3192 (N10760, N10707, N10553);
  or OR2_3193 (N10761, N10708, N10554);
  or OR2_3194 (N10762, N10709, N10555);
  or OR2_3195 (N10763, N10710, N10556);
  or OR2_3209 (N10837, N10730, N10587);
  or OR2_3210 (N10839, N10731, N10588);
  or OR2_3277 (N10905, N10864, N10765);
  or OR2_3278 (N10906, N10865, N10766);
  or OR2_3279 (N10907, N10866, N10767);
  or OR2_3280 (N10908, N10867, N10768);
  or OR2_3485 (N11299, N11288, N11278);
  or OR2_3486 (N11302, N11289, N11280);
  or OR2_3495 (N11317, N11309, N11298);
  or OR2_3498 (N11323, N11308, N11316);
  or OR3_922 (N4303, N1167, N2866, N3122);
  or OR3_2044 (N8204, N3173, N6844, N6865);
  or OR3_2420 (N9107, N4549, N8345, N8346);
  or OR3_2430 (N9169, N4661, N8441, N8442);
  or OR3_2646 (N9632, N4570, N8357, N9287);
  or OR3_2893 (N10119, N9791, N10042, N10043);
  or OR3_2907 (N10148, N9791, N10060, N10061);
  or OR3_3026 (N10412, N3195, N6864, N10289);
  or OR3_3030 (N10425, N3107, N6782, N10280);
  or OR3_3136 (N10665, N4682, N8456, N10596);
  or OR4_2019 (N7649, N3168, N6836, N6837, N6838);
  or OR4_2027 (N7825, N3361, N7060, N7061, N7062);
  or OR4_2030 (N8114, N3101, N6777, N6778, N6779);
  or OR4_2036 (N8146, N3169, N6839, N6840, N6841);
  or OR4_2038 (N8166, N3189, N6859, N6860, N6861);
  or OR4_2371 (N8898, N4544, N8337, N8338, N8339);
  or OR4_2378 (N8950, N4630, N8409, N8410, N8411);
  or OR4_2382 (N8963, N4656, N8433, N8434, N8435);
  or OR4_2392 (N9029, N4756, N8545, N8546, N8547);
  or OR4_2418 (N9099, N4545, N8340, N8341, N8342);
  or OR4_2428 (N9161, N4657, N8436, N8437, N8438);
  or OR4_2438 (N9203, N4678, N8454, N8455, N8513);
  or OR4_2645 (N9629, N4566, N8355, N8356, N9286);
  or OR4_2667 (N9679, N4566, N8355, N8356, N9315);
  or OR4_2892 (N10116, N9265, N10039, N10040, N10041);
  or OR4_2905 (N10140, N8943, N10055, N10056, N9790);
  or OR4_2906 (N10141, N9265, N10057, N10058, N10059);
  or OR4_3025 (N10409, N3189, N6859, N6860, N10288);
  or OR4_3029 (N10422, N3101, N6777, N6778, N10279);
  or OR4_3135 (N10662, N4678, N8454, N8455, N10595);
  or OR4_3183 (N10739, N10648, N10649, N10581, N10582);
  or OR4_3421 (N11205, N11152, N11153, N11154, N11155);
  or OR4_3452 (N11252, N11222, N11223, N11224, N11225);
  or OR4_3453 (N11257, N11226, N11227, N11228, N11229);
  or g1 (n_316, N3126, N8818);
  or g2 (n_317, N9732, N10013);
  or g3 (N10101, N10014, N10015, n_316, n_317);
  and g4 (n_318, N367, N9754);
  and g5 (N10015, N9344, N8307, N8269, n_318);
  or g6 (n_319, N3096, N6766);
  or g7 (N7609, N6767, N6768, N6769, n_319);
  and g8 (n_320, N5670, N5654);
  and g9 (N6769, N5632, N3114, N5640, n_320);
  and g10 (n_321, N5640, N5683);
  and g11 (N6784, N5654, N5632, N5670, n_321);
  and g12 (n_322, N5807, N5856);
  and g13 (N6881, N5821, N5799, N5837, n_322);
  and g14 (n_323, N7149, N7180);
  and g15 (N8444, N7159, N7142, N7170, n_323);
  and g16 (n_324, N6936, N8326);
  and g17 (N9280, N6946, N6929, N6957, n_324);
  or g18 (n_325, N3184, N6848);
  or g19 (N7655, N6849, N6850, N6851, n_325);
  or g20 (n_326, N4674, N8447);
  or g21 (N8966, N8448, N8449, N8450, n_326);
  or g22 (n_327, N4562, N8348);
  or g23 (N8902, N8349, N8350, N8351, n_327);
  and g24 (n_328, N5837, N5821);
  and g25 (N6851, N5799, N3202, N5807, n_328);
  and g26 (n_329, N7170, N7159);
  and g27 (N8450, N7142, N4687, N7149, n_329);
  and g28 (n_330, N6957, N6946);
  and g29 (N8351, N6929, N5960, N6936, n_330);
  or g30 (n_331, N4193, N8960);
  or g31 (n_332, N9526, N10016);
  or g32 (N10102, N10017, N9734, n_331, n_332);
  and g33 (n_333, N89, N9408);
  and g34 (N9734, N9332, N8394, N8421, n_333);
  or g35 (n_334, N3370, N7103);
  or g36 (N7852, N7104, N7105, N7106, n_334);
  and g37 (n_335, N7057, N6022);
  and g39 (N8394, N6009, N6003, n_335, n_336);
  and g40 (N7104, N6047, N6041, N2662, N2450);
  and g41 (n_337, N6056, N6052);
  and g42 (n_338, N6041, N2654);
  and g43 (N7106, N628, N6047, n_337, n_338);
  and g44 (N7061, N5996, N5991, N2753, N2470);
  and g45 (n_339, N6059, N6056);
  and g46 (N7100, N6052, N6047, N6041, n_339);
  and g47 (n_340, N7099, N7095);
  and g48 (N8412, N7091, N7086, N7080, n_340);
  and g49 (n_341, N7377, N7373);
  and g50 (N8548, N7369, N7364, N7358, n_341);
  or g51 (n_342, N3365, N7064);
  or g52 (N7826, N7065, N7066, N7067, n_342);
  and g53 (N8410, N7073, N7068, N3440, N2696);
  or g54 (n_343, N4637, N8415);
  or g55 (N8956, N8416, N8417, N8418, n_343);
  and g56 (N8546, N7351, N7346, N3474, N3255);
  or g57 (n_344, N4760, N8551);
  or g58 (N9035, N8552, N8553, N8554, n_344);
  and g59 (N7065, N6009, N6003, N2737, N2546);
  and g60 (n_336, N6018, N6014);
  and g61 (n_346, N6003, N2729);
  and g62 (N7067, N2538, N6009, n_336, n_346);
  and g63 (N8416, N7086, N7080, N3424, N3307);
  and g64 (n_347, N7095, N7091);
  and g65 (n_348, N7080, N3416);
  and g66 (N8418, N3299, N7086, n_347, n_348);
  and g67 (N8552, N7364, N7358, N3458, N2611);
  and g68 (n_349, N7373, N7369);
  and g69 (n_350, N7358, N2680);
  and g70 (N8554, N3381, N7364, n_349, n_350);
  or g72 (n_352, N9736, N10020);
  or g73 (N10104, N10021, N10022, n_316, n_352);
  and g74 (n_353, N367, N9775);
  and g75 (N10022, N9385, N8298, N8262, n_353);
  and g77 (N6762, N5654, N5640, N5632, N6783);
  and g79 (N6845, N5821, N5807, N5799, N6866);
  and g81 (N8497, N7159, N7149, N7142, N8518);
  and g83 (N9307, N6946, N6936, N6929, N9318);
  or g84 (n_358, N4563, N8352);
  or g85 (N9626, N8353, N8354, N9285, n_358);
  and g87 (N9285, N6946, N6957, N6936, N9288);
  or g89 (N10406, N6853, N6854, N10287, n_360);
  and g91 (N10287, N5821, N5837, N5807, N10290);
  or g93 (N10419, N6771, N6772, N10278, n_362);
  and g95 (N10278, N5654, N5670, N5640, N10281);
  or g97 (N10659, N8452, N8453, N10594, n_364);
  and g99 (N10594, N7159, N7170, N7149, N10597);
  or g100 (n_360, N3185, N6852);
  or g101 (N8169, N6853, N6854, N6855, n_360);
  or g102 (n_362, N3097, N6770);
  or g103 (N8117, N6771, N6772, N6773, n_362);
  or g104 (n_364, N4675, N8451);
  or g105 (N9206, N8452, N8453, N8507, n_364);
  or g107 (N9685, N8353, N8354, N9314, n_358);
endmodule

